

module Cache #(
   parameter CPU_WIDTH = 32,

)(
    
);

endmodule //Cache
