module div (
    
);

endmodule //div