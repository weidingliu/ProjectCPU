`define RestEn 1'b1
`define RestDis 1'b0
`define false 1'b0
`define true 1'b1
`define ctrl_width 186
`define ex_ctrl_width 213
`define mem_ctrl_width 103