`define RestEn 1'b1
`define RestDis 1'b0
`define ctrl_width 166