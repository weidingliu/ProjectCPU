module mul (
    ports
);
    
endmodule