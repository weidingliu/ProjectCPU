/*
* this is booth-2 multiplier,use chisel to convert verilog,here is verilog code
*
*/

module Partial_product(
  input  [2:0]  io_y_3,
  input  [67:0] io_x,
  output [67:0] io_p,
  output        io_c
);
  wire  _io_p_T = io_y_3 == 3'h0; // @[MUL.scala 26:13]
  wire  _io_p_T_1 = io_y_3 == 3'h1; // @[MUL.scala 27:13]
  wire  _io_p_T_2 = io_y_3 == 3'h2; // @[MUL.scala 28:13]
  wire  _io_p_T_3 = io_y_3 == 3'h3; // @[MUL.scala 29:13]
  wire [68:0] _io_p_T_4 = {io_x, 1'h0}; // @[MUL.scala 29:36]
  wire  _io_p_T_5 = io_y_3 == 3'h4; // @[MUL.scala 30:13]
  wire [68:0] _io_p_T_7 = ~_io_p_T_4; // @[MUL.scala 30:31]
  wire  _io_p_T_8 = io_y_3 == 3'h5; // @[MUL.scala 31:13]
  wire [67:0] _io_p_T_9 = ~io_x; // @[MUL.scala 31:32]
  wire  _io_p_T_10 = io_y_3 == 3'h6; // @[MUL.scala 32:13]
  wire [67:0] _io_p_T_14 = _io_p_T_10 ? _io_p_T_9 : 68'h0; // @[Mux.scala 101:16]
  wire [67:0] _io_p_T_15 = _io_p_T_8 ? _io_p_T_9 : _io_p_T_14; // @[Mux.scala 101:16]
  wire [68:0] _io_p_T_16 = _io_p_T_5 ? _io_p_T_7 : {{1'd0}, _io_p_T_15}; // @[Mux.scala 101:16]
  wire [68:0] _io_p_T_17 = _io_p_T_3 ? _io_p_T_4 : _io_p_T_16; // @[Mux.scala 101:16]
  wire [68:0] _io_p_T_18 = _io_p_T_2 ? {{1'd0}, io_x} : _io_p_T_17; // @[Mux.scala 101:16]
  wire [68:0] _io_p_T_19 = _io_p_T_1 ? {{1'd0}, io_x} : _io_p_T_18; // @[Mux.scala 101:16]
  wire [68:0] _io_p_T_20 = _io_p_T ? 69'h0 : _io_p_T_19; // @[Mux.scala 101:16]
  wire  _io_c_T_12 = _io_p_T_3 ? 1'h0 : _io_p_T_5 | (_io_p_T_8 | _io_p_T_10); // @[Mux.scala 101:16]
  wire  _io_c_T_13 = _io_p_T_2 ? 1'h0 : _io_c_T_12; // @[Mux.scala 101:16]
  wire  _io_c_T_14 = _io_p_T_1 ? 1'h0 : _io_c_T_13; // @[Mux.scala 101:16]
  assign io_p = _io_p_T_20[67:0]; // @[MUL.scala 25:8]
  assign io_c = _io_p_T ? 1'h0 : _io_c_T_14; // @[Mux.scala 101:16]
endmodule
module Booth_MUL(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_ctrl_flow_flush,
  input         io_in_bits_ctrl_flow_mulw,
  input  [1:0]  io_in_bits_ctrl_flow_mul_sign,
  input  [31:0] io_in_bits_ctrl_data_src1,
  input  [31:0] io_in_bits_ctrl_data_src2,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result_result_hi,
  output [31:0] io_out_bits_result_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] partial_io_y_3; // @[MUL.scala 134:23]
  wire [67:0] partial_io_x; // @[MUL.scala 134:23]
  wire [67:0] partial_io_p; // @[MUL.scala 134:23]
  wire  partial_io_c; // @[MUL.scala 134:23]
  reg [33:0] multiplier; // @[MUL.scala 130:27]
  reg [67:0] multiplicand; // @[MUL.scala 131:29]
  reg [67:0] p; // @[MUL.scala 132:18]
  reg [5:0] count; // @[MUL.scala 133:22]
  wire  sign = io_in_bits_ctrl_data_src1[31]; // @[util.scala 10:19]
  wire [32:0] _T = {sign,io_in_bits_ctrl_data_src1}; // @[Cat.scala 33:92]
  wire  sign_1 = io_in_bits_ctrl_data_src2[31]; // @[util.scala 10:19]
  wire [32:0] _T_1 = {sign_1,io_in_bits_ctrl_data_src2}; // @[Cat.scala 33:92]
  wire [32:0] _T_3 = {1'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 33:92]
  wire [32:0] _T_4 = {1'h0,io_in_bits_ctrl_data_src1}; // @[Cat.scala 33:92]
  wire  _src1_T = 2'h0 == io_in_bits_ctrl_flow_mul_sign; // @[util.scala 31:32]
  wire  _src1_T_1 = 2'h1 == io_in_bits_ctrl_flow_mul_sign; // @[util.scala 31:32]
  wire  _src1_T_2 = 2'h3 == io_in_bits_ctrl_flow_mul_sign; // @[util.scala 31:32]
  wire [32:0] _src1_T_3 = _src1_T ? _T : 33'h0; // @[Mux.scala 27:73]
  wire [32:0] _src1_T_4 = _src1_T_1 ? _T : 33'h0; // @[Mux.scala 27:73]
  wire [32:0] _src1_T_5 = _src1_T_2 ? _T_4 : 33'h0; // @[Mux.scala 27:73]
  wire [32:0] _src1_T_6 = _src1_T_3 | _src1_T_4; // @[Mux.scala 27:73]
  wire [32:0] src1 = _src1_T_6 | _src1_T_5; // @[Mux.scala 27:73]
  wire [32:0] _src2_T_3 = _src1_T ? _T_1 : 33'h0; // @[Mux.scala 27:73]
  wire [32:0] _src2_T_4 = _src1_T_1 ? _T_3 : 33'h0; // @[Mux.scala 27:73]
  wire [32:0] _src2_T_5 = _src1_T_2 ? _T_3 : 33'h0; // @[Mux.scala 27:73]
  wire [32:0] _src2_T_6 = _src2_T_3 | _src2_T_4; // @[Mux.scala 27:73]
  wire [32:0] src2 = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  wire  _count_T_1 = ~io_in_bits_ctrl_flow_flush & io_in_valid; // @[MUL.scala 146:44]
  wire [5:0] _count_T_5 = count + 6'h2; // @[MUL.scala 146:81]
  wire [33:0] _multiplier_T = {src2,1'h0}; // @[Cat.scala 33:92]
  wire [67:0] _multiplicand_T_1 = {1'h0,src1,34'h0}; // @[Cat.scala 33:92]
  wire [67:0] _temp_T_1 = p + partial_io_p; // @[MUL.scala 154:18]
  wire [67:0] _GEN_6 = {{67'd0}, partial_io_c}; // @[MUL.scala 154:28]
  wire [67:0] temp = _temp_T_1 + _GEN_6; // @[MUL.scala 154:28]
  wire  p_sign = temp[67]; // @[util.scala 10:19]
  wire [1:0] _p_T_2 = p_sign ? 2'h3 : 2'h0; // @[Bitwise.scala 77:12]
  wire [67:0] _p_T_3 = {_p_T_2,temp[67:2]}; // @[Cat.scala 33:92]
  Partial_product partial ( // @[MUL.scala 134:23]
    .io_y_3(partial_io_y_3),
    .io_x(partial_io_x),
    .io_p(partial_io_p),
    .io_c(partial_io_c)
  );
  assign io_in_ready = 1'h1; // @[MUL.scala 164:15]
  assign io_out_valid = count == 6'h24 & io_in_bits_ctrl_flow_mulw | count == 6'h24; // @[MUL.scala 163:84]
  assign io_out_bits_result_result_hi = p[63:32]; // @[MUL.scala 165:36]
  assign io_out_bits_result_result_lo = p[31:0]; // @[MUL.scala 166:36]
  assign partial_io_y_3 = multiplier[2:0]; // @[MUL.scala 160:31]
  assign partial_io_x = multiplicand; // @[MUL.scala 161:16]
  always @(posedge clock) begin
    if (reset) begin // @[MUL.scala 130:27]
      multiplier <= 34'h0; // @[MUL.scala 130:27]
    end else if (_count_T_1) begin // @[MUL.scala 147:51]
      if (count == 6'h0) begin // @[MUL.scala 148:25]
        multiplier <= _multiplier_T; // @[MUL.scala 149:18]
      end else begin
        multiplier <= {{2'd0}, multiplier[33:2]}; // @[MUL.scala 156:18]
      end
    end
    if (reset) begin // @[MUL.scala 131:29]
      multiplicand <= 68'h0; // @[MUL.scala 131:29]
    end else if (_count_T_1) begin // @[MUL.scala 147:51]
      if (count == 6'h0) begin // @[MUL.scala 148:25]
        multiplicand <= _multiplicand_T_1; // @[MUL.scala 150:20]
      end
    end
    if (reset) begin // @[MUL.scala 132:18]
      p <= 68'h0; // @[MUL.scala 132:18]
    end else if (_count_T_1) begin // @[MUL.scala 147:51]
      if (count == 6'h0) begin // @[MUL.scala 148:25]
        p <= 68'h0; // @[MUL.scala 151:9]
      end else begin
        p <= _p_T_3; // @[MUL.scala 155:9]
      end
    end
    if (reset) begin // @[MUL.scala 133:22]
      count <= 6'h0; // @[MUL.scala 133:22]
    end else if (~io_in_bits_ctrl_flow_flush & io_in_valid & ~io_out_valid) begin // @[MUL.scala 146:15]
      count <= _count_T_5;
    end else begin
      count <= 6'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  multiplier = _RAND_0[33:0];
  _RAND_1 = {3{`RANDOM}};
  multiplicand = _RAND_1[67:0];
  _RAND_2 = {3{`RANDOM}};
  p = _RAND_2[67:0];
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule



// ###############################################################################################################3

/*then is scala code*/

// import chisel3._
// import chisel3.util._

// object Siganle{
//   val ss = "b00".U
//   val su = "b01".U
//   val uu = "b11".U
// }

// class Partial_product (booth_bit : Int = 3, mul_len: Int)extends Module{
//   val io = IO(new Bundle() {
//     val y_3 = Input(UInt(booth_bit.W))
//     val x = Input(UInt(((mul_len+2)*2).W))
//     val p = Output(UInt(((mul_len+2)*2).W))
//     val c = Output(UInt(1.W))
//   })


//   io.p := MuxCase(0.U(((mul_len+2)*2).W),Seq(
//     (io.y_3 === "b000".U) -> 0.U(((mul_len+2)*2).W),
//     (io.y_3 === "b001".U) -> io.x,
//     (io.y_3 === "b010".U) -> io.x,
//     (io.y_3 === "b011".U) -> (io.x << 1),
//     (io.y_3 === "b100".U) -> (~(io.x << 1)),
//     (io.y_3 === "b101".U) -> ((~io.x)),
//     (io.y_3 === "b110".U) -> (~io.x),
//     (io.y_3 === "b111".U) -> 0.U(((mul_len+2)*2).W),

//   ))
//   io.c := MuxCase(0.U(1.W), Seq(
//     (io.y_3 === "b000".U) -> 0.U(1.W),
//     (io.y_3 === "b001".U) -> 0.U(1.W),
//     (io.y_3 === "b010".U) -> 0.U(1.W),
//     (io.y_3 === "b011".U) -> 0.U(1.W),
//     (io.y_3 === "b100".U) -> 1.U(1.W),
//     (io.y_3 === "b101".U) -> 1.U(1.W),
//     (io.y_3 === "b110".U) -> 1.U(1.W),
//     (io.y_3 === "b111".U) -> 0.U(1.W),

//   ))
// }
// object Partial_product{
//     def apply(booth_bit : Int = 3, mul_len: Int,y_3:UInt,x:UInt) ={
//       val m = Module(new Partial_product(booth_bit,mul_len))
//       m.io.y_3 := y_3
//       m.io.x := x
//       (m.io.p,m.io.c)
//     }
// }

// class Booth_MUL(booth_bit : Int = 3, mul_len: Int) extends Module{
//   val io = IO(new Bundle() {
//     val in = Flipped(Decoupled(new MUL_IN(mul_len)))
//     val out = Decoupled(new MUL_OUT(mul_len))
//   })

//   val multiplier = RegInit(0.U(((mul_len+2)).W))
//   val multiplicand = RegInit(0.U(((mul_len+2)*2).W))
//   val p = RegInit(0.U(((mul_len+2)*2).W))
//   val count = RegInit(0.U(log2Ceil(mul_len+4).W))
//   val partial = Module(new Partial_product(booth_bit = 3,mul_len=mul_len))
//   val partial_c = partial.io.c
//   val partial_p = partial.io.p

//   val list_table = List(
//     (Siganle.ss) -> (SIgEXtend(io.in.bits.ctrl_data.src1,mul_len+1),SIgEXtend(io.in.bits.ctrl_data.src2,mul_len+1)),
//     (Siganle.su) -> (SIgEXtend(io.in.bits.ctrl_data.src1,mul_len+1),ZeroEXtend(io.in.bits.ctrl_data.src2,mul_len+1)),
//     (Siganle.uu) -> (ZeroEXtend(io.in.bits.ctrl_data.src1,mul_len+1),ZeroEXtend(io.in.bits.ctrl_data.src2,mul_len+1)),
//   )
//   val src1 = LookupTree(io.in.bits.ctrl_flow.mul_sign,list_table.map(p => (p._1,p._2._1)))
//   val src2 = LookupTree(io.in.bits.ctrl_flow.mul_sign,list_table.map(p => (p._1,p._2._2)))

  
  // count := Mux(!io.in.bits.ctrl_flow.flush && io.in.valid && !io.out.valid,count+2.U,0.U)
  // when(!io.in.bits.ctrl_flow.flush && io.in.valid){
  //   when (count === 0.U){
  //     multiplier := Cat(src2, Fill(1, 0.U))//xlen+2
  //     multiplicand := Cat(Fill(1,0.U),src1, Fill(mul_len + 2, 0.U))
  //     p := 0.U
  //   }
  //   .otherwise {
  //     val temp =p+partial_p+partial_c
  //     p := SIgEXtend(temp((mul_len+2)*2-1,2),(mul_len+2)*2)
  //     multiplier := multiplier >> 2
  //   }
  // }

  // partial.io.y_3 := multiplier(2,0)
  // partial.io.x := multiplicand

  // io.out.valid := Mux((count === ((mul_len+2) + 2).U && io.in.bits.ctrl_flow.mulw) || count === ((mul_len+2) + 2).U, true.B, false.B)
  // io.in.ready := true.B
  // io.out.bits.result.result_hi := p(mul_len * 2 -1, mul_len)
  // io.out.bits.result.result_lo := p(mul_len -1 , 0)

// }


// ############################### here is walloc_booth mul ################################################

// class Improved_Partial_product(mul_len : Int)extends Module{
//   val io = IO(new Bundle(){
//     val y_3 = Input(UInt(3.W))
//     val x = Input(UInt((mul_len+2).W))
//     val p = Output(UInt((mul_len+2).W))
//     val carry = Output(UInt(2.W))
// })
//   io.p := MuxCase(0.U((mul_len + 2).W), Seq(
//     (io.y_3 === "b000".U) -> 0.U(((mul_len + 2)).W),
//     (io.y_3 === "b001".U) -> io.x,
//     (io.y_3 === "b010".U) -> io.x,
//     (io.y_3 === "b011".U) -> (io.x << 1),
//     (io.y_3 === "b100".U) -> ((~io.x) << 1),
//     (io.y_3 === "b101".U) -> (~io.x),
//     (io.y_3 === "b110".U) -> (~io.x),
//     (io.y_3 === "b111".U) -> 0.U(((mul_len + 2)).W),

//   ))
//   io.carry := MuxCase(0.U(2.W), Seq(
//     (io.y_3 === "b000".U) -> "b00".U(2.W),
//     (io.y_3 === "b001".U) -> "b00".U(2.W),
//     (io.y_3 === "b010".U) -> "b00".U(2.W),
//     (io.y_3 === "b011".U) -> "b00".U(2.W),
//     (io.y_3 === "b100".U) -> "b10".U(2.W),
//     (io.y_3 === "b101".U) -> "b01".U(2.W),
//     (io.y_3 === "b110".U) -> "b01".U(2.W),
//     (io.y_3 === "b111".U) -> "b00".U(2.W),
//   ))
// }
// object Improved_Partial_product{
//     def apply( mul_len: Int,y_3:UInt,x:UInt) ={
//       val m = Module(new Improved_Partial_product(mul_len))
//       m.io.y_3 := y_3
//       m.io.x := x
//       (m.io.p,m.io.carry)
//     }
// }

// class Adder extends Module with Paramete{
//   val io = IO(new Bundle() {
//     val x1 = Input(UInt(1.W))
//     val x2 = Input(UInt(1.W))
//     val x3 = Input(UInt(1.W))
//     val s = Output(UInt(1.W))
//     val cout = Output(UInt(1.W))
//   })
//   io.s := io.x1 ^ io.x2 ^ io.x3
//   io.cout := (io.x1 & io.x2) | (io.x1 & io.x3) | (io.x2 & io.x3)
// }

// object Adder  {
//   def apply(x1:UInt,x2:UInt,x3:UInt) ={
//     val m = Module(new Adder)
//     m.io.x1 := x1
//     m.io.x2 := x2
//     m.io.x3 := x3
// //    Cat(m.io.s,m.io.c)
//     (m.io.s,m.io.cout)

// //    s := m.io.s
// //    c := m.io.c
//   }
// }

// class Half_Adder extends Module{
//   val io = IO(new Bundle() {
//     val in = Input(Vec(2,Bool()))
//     val out = Output(Vec(2,Bool()))
//   })
//   io.out(0) := io.in(0) ^ io.in(1)
//   io.out(1) := io.in(0) & io.in(1)
// }
// object Half_Adder{
//   def apply(in1:Bool,in2:Bool): (Bool,Bool) = {
//     val m = Module(new Half_Adder)
//     m.io.in(0) := in1
//     m.io.in(1) := in2
//     (m.io.out(0) ,m.io.out(1))
//   }
// }

// class Booth_Walloc_MUL (mul_len:Int) extends Module with Paramete{
//   val io = IO(new Bundle() {
//     val in = Flipped(Decoupled(new MUL_IN(mul_len)))
//     val out = Decoupled(new MUL_OUT(mul_len))
//   })
//   def max_col (y:Array[Seq[Bool]]): Int = {
//     var max_size = 0
//     for(i <- 0 until y.size){
//       if(max_size < y(i).size) max_size = y(i).size
//     }
//     max_size
//   }
//   def array_take(y:Seq[Bool],x:Seq[Bool]): Seq[Bool] ={
//     if(y == null){
//       x
//     }
//     else{
//       y ++ x
//     }
//   }
//   def select_elem(x:Array[Seq[Bool]],index:Int): Seq[Bool]={
//     var temp = Seq[Bool]()
//     for(i <- 0 until x.size){
//       temp = temp :+ x(i)(index)
//     }
// //    Cat(temp.reverse)
//     temp
//   }

//   def Add_Onecolmn(col:Seq[Bool],cin:Seq[Bool]): (Seq[Bool],Seq[Bool]) = {
//     var sum = Seq[Bool]()
//     var cout = Seq[Bool]()

//     col.size match {
//       case 1 => {
//         sum = col ++ cin
//       }
//       case 2 => {
//         val (s,c) = Half_Adder(col(0),col(1))
//         sum = Seq(s) ++ cin
//         cout = Seq(c)
//       }
//       case 3 => {
//         val (s,c) = Adder(col(0),col(1),col(2))
//         sum = Seq(s.asBool) ++ cin
//         cout = Seq(c.asBool)
//       }
//       case n => {
//         val count_1 = if(cin.nonEmpty) Seq(cin.head) else Nil
//         val count_2 = if(cin.nonEmpty) cin.drop(1) else Nil
//         val (s_1,c_1) = Add_Onecolmn(col take 3,count_1)
//         val (s_2,c_2) = Add_Onecolmn(col drop 3,count_2)
//         sum = s_1 ++ s_2
//         cout = c_1 ++ c_2
//       }
//     }
//     (sum,cout)
//   }
//   def Add_All(cols: Array[Seq[Bool]],depth:Int): (UInt,UInt) ={

//     if(max_col(cols) <= 2){
//       val sum = Cat(select_elem(cols,0).reverse)
//       var k = 0
//       while(cols(k).size == 1) k = k+1
//       val carry = Cat(select_elem(cols.drop(k),1).reverse)
// //      println(depth)
//       (sum,Cat(carry,Fill(k,0.U(1.W))))
//     }
//     else {
//       val columns_next = Array.fill(cols.size)(Seq[Bool]())
//       var cout = Seq[Bool]()
//       for(i<-0 until cols.size){
//         val (s,c) = Add_Onecolmn(cols(i),cout)
//         columns_next(i) = s
//         cout = c
//       }
// //      println(depth)
//       val next_layer = if(depth == 3) columns_next.map(col => col.map(x => RegEnable(x,io.in.valid))) else columns_next
//       Add_All(next_layer,depth+1)
//     }
//   }

//   // src2 is Double sign bit
//   val list_table = List(
//     (Siganle.ss) -> (Cat(SIgEXtend(io.in.bits.ctrl_data.src1, mul_len + 2),Fill(1,0.U)), SIgEXtend(io.in.bits.ctrl_data.src2, mul_len + 2)),
//     (Siganle.su) -> (Cat(SIgEXtend(io.in.bits.ctrl_data.src1, mul_len + 2),Fill(1,0.U)), ZeroEXtend(io.in.bits.ctrl_data.src2, mul_len + 2)),
//     (Siganle.uu) -> (Cat(ZeroEXtend(io.in.bits.ctrl_data.src1, mul_len + 2),Fill(1,0.U)), ZeroEXtend(io.in.bits.ctrl_data.src2, mul_len + 2)),
//   )
//   val src1 = LookupTree(io.in.bits.ctrl_flow.mul_sign, list_table.map(p => (p._1, p._2._1)))
//   val src2 = LookupTree(io.in.bits.ctrl_flow.mul_sign, list_table.map(p => (p._1, p._2._2)))

//   val partial_product_array = new Array[Seq[Bool]]((mul_len +2 )*2-1)
// //  val last_c = Seq[UInt]
//   var next_c = 0.U(2.W)
//   for (i<-0 until (mul_len+2) by 2){
//     val (p,c_p) = Improved_Partial_product(mul_len,src1(i+2,i),src2)
//     for(j<-0 until (mul_len+2)){
//       partial_product_array(j + i) = array_take(partial_product_array(j + i) , Seq(p(j)))
//       if(j == mul_len +1 && i != 0 && i != mul_len){
//         partial_product_array(j + i +1) = array_take(partial_product_array(j + i +1) , Seq(!p(j)))
//         partial_product_array(j + i +2) = array_take(partial_product_array(j + i +2) , Seq(1.B))
//       }
//       if(j == mul_len +1 && i == 0){
//         partial_product_array(j + i + 1) = array_take(partial_product_array(j + i + 1), Seq(p(j)))
//         partial_product_array(j + i + 2) = array_take(partial_product_array(j + i + 2), Seq(p(j)))
//         partial_product_array(j + i + 3) = array_take(partial_product_array(j + i + 3), Seq(!p(j)))
//       }
//       if(j == mul_len +1 && i == mul_len){
//         partial_product_array(j + i +1) = array_take(partial_product_array(j + i +1) , Seq(!p(j)))
//       }
//     }
//     if (i != 0) {
//       partial_product_array(i - 1) = array_take(partial_product_array(i - 1), Seq(next_c(1)))
//       partial_product_array(i - 2) = array_take(partial_product_array(i - 2), Seq(next_c(0)))
//     }
//     next_c = c_p
//   }
// //for(i<-0 until partial_product_array.size){
// //  println(i.toString +" "+ partial_product_array(i).size.toString)
// //}
// //  println(partial_product_array.size)
//   val cols_reg = partial_product_array.map(col => col.map(x => RegEnable(x,io.in.valid)))
//   val (sum,cout) = Add_All(cols_reg,0)

//   val result = sum + cout

//   val count = RegInit(0.U(8.W))
//   val s = count === 2.U(8.W)
//   count := Mux(!io.in.bits.ctrl_flow.flush && io.in.valid && !io.out.valid,count+1.U,0.U)
// //  when(io.in.valid){
// //    count := count +1.U(8.W)
// //  }.otherwise{
// //    count := 0.U(8.W)
// //  }

//   io.out.bits.result.result_hi := result(mul_len * 2-1,mul_len)
//   io.out.bits.result.result_lo:= result(mul_len -1,0)
//   io.out.valid := Mux(s,true.B,false.B)
//   io.in.ready := true.B
// }


module Improved_Partial_product(
  input  [2:0]  io_y_3,
  input  [33:0] io_x,
  output [33:0] io_p,
  output [1:0]  io_carry
);
  wire  _io_p_T = io_y_3 == 3'h0; // @[MUL.scala 58:13]
  wire  _io_p_T_1 = io_y_3 == 3'h1; // @[MUL.scala 59:13]
  wire  _io_p_T_2 = io_y_3 == 3'h2; // @[MUL.scala 60:13]
  wire  _io_p_T_3 = io_y_3 == 3'h3; // @[MUL.scala 61:13]
  wire [34:0] _io_p_T_4 = {io_x, 1'h0}; // @[MUL.scala 61:36]
  wire  _io_p_T_5 = io_y_3 == 3'h4; // @[MUL.scala 62:13]
  wire [33:0] _io_p_T_6 = ~io_x; // @[MUL.scala 62:32]
  wire [34:0] _io_p_T_7 = {_io_p_T_6, 1'h0}; // @[MUL.scala 62:39]
  wire  _io_p_T_8 = io_y_3 == 3'h5; // @[MUL.scala 63:13]
  wire  _io_p_T_10 = io_y_3 == 3'h6; // @[MUL.scala 64:13]
  wire [33:0] _io_p_T_14 = _io_p_T_10 ? _io_p_T_6 : 34'h0; // @[Mux.scala 101:16]
  wire [33:0] _io_p_T_15 = _io_p_T_8 ? _io_p_T_6 : _io_p_T_14; // @[Mux.scala 101:16]
  wire [34:0] _io_p_T_16 = _io_p_T_5 ? _io_p_T_7 : {{1'd0}, _io_p_T_15}; // @[Mux.scala 101:16]
  wire [34:0] _io_p_T_17 = _io_p_T_3 ? _io_p_T_4 : _io_p_T_16; // @[Mux.scala 101:16]
  wire [34:0] _io_p_T_18 = _io_p_T_2 ? {{1'd0}, io_x} : _io_p_T_17; // @[Mux.scala 101:16]
  wire [34:0] _io_p_T_19 = _io_p_T_1 ? {{1'd0}, io_x} : _io_p_T_18; // @[Mux.scala 101:16]
  wire [34:0] _io_p_T_20 = _io_p_T ? 35'h0 : _io_p_T_19; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_9 = _io_p_T_10 ? 2'h1 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_10 = _io_p_T_8 ? 2'h1 : _io_carry_T_9; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_11 = _io_p_T_5 ? 2'h2 : _io_carry_T_10; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_12 = _io_p_T_3 ? 2'h0 : _io_carry_T_11; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_13 = _io_p_T_2 ? 2'h0 : _io_carry_T_12; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_14 = _io_p_T_1 ? 2'h0 : _io_carry_T_13; // @[Mux.scala 101:16]
  assign io_p = _io_p_T_20[33:0]; // @[MUL.scala 57:8]
  assign io_carry = _io_p_T ? 2'h0 : _io_carry_T_14; // @[Mux.scala 101:16]
endmodule
module Half_Adder(
  input   io_in_0,
  input   io_in_1,
  output  io_out_0,
  output  io_out_1
);
  assign io_out_0 = io_in_0 ^ io_in_1; // @[MUL.scala 119:25]
  assign io_out_1 = io_in_0 & io_in_1; // @[MUL.scala 120:25]
endmodule
module Adder(
  input   io_x1,
  input   io_x2,
  input   io_x3,
  output  io_s,
  output  io_cout
);
  assign io_s = io_x1 ^ io_x2 ^ io_x3; // @[MUL.scala 96:25]
  assign io_cout = io_x1 & io_x2 | io_x1 & io_x3 | io_x2 & io_x3; // @[MUL.scala 97:48]
endmodule
module Booth_Walloc_MUL(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_ctrl_flow_flush,
  input         io_in_bits_ctrl_flow_mulw,
  input  [1:0]  io_in_bits_ctrl_flow_mul_sign,
  input  [31:0] io_in_bits_ctrl_data_src1,
  input  [31:0] io_in_bits_ctrl_data_src2,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_result_result_hi,
  output [31:0] io_out_bits_result_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] m_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_1_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_1_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_1_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_1_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_2_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_2_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_2_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_2_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_3_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_3_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_3_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_3_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_4_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_4_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_4_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_4_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_5_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_5_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_5_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_5_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_6_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_6_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_6_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_6_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_7_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_7_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_7_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_7_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_8_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_8_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_8_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_8_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_9_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_9_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_9_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_9_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_10_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_10_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_10_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_10_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_11_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_11_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_11_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_11_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_12_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_12_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_12_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_12_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_13_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_13_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_13_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_13_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_14_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_14_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_14_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_14_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_15_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_15_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_15_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_15_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_16_io_y_3; // @[MUL.scala 81:21]
  wire [33:0] m_16_io_x; // @[MUL.scala 81:21]
  wire [33:0] m_16_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_16_io_carry; // @[MUL.scala 81:21]
  wire  m_17_io_in_0; // @[MUL.scala 124:19]
  wire  m_17_io_in_1; // @[MUL.scala 124:19]
  wire  m_17_io_out_0; // @[MUL.scala 124:19]
  wire  m_17_io_out_1; // @[MUL.scala 124:19]
  wire  m_18_io_in_0; // @[MUL.scala 124:19]
  wire  m_18_io_in_1; // @[MUL.scala 124:19]
  wire  m_18_io_out_0; // @[MUL.scala 124:19]
  wire  m_18_io_out_1; // @[MUL.scala 124:19]
  wire  m_19_io_x1; // @[MUL.scala 102:19]
  wire  m_19_io_x2; // @[MUL.scala 102:19]
  wire  m_19_io_x3; // @[MUL.scala 102:19]
  wire  m_19_io_s; // @[MUL.scala 102:19]
  wire  m_19_io_cout; // @[MUL.scala 102:19]
  wire  m_20_io_x1; // @[MUL.scala 102:19]
  wire  m_20_io_x2; // @[MUL.scala 102:19]
  wire  m_20_io_x3; // @[MUL.scala 102:19]
  wire  m_20_io_s; // @[MUL.scala 102:19]
  wire  m_20_io_cout; // @[MUL.scala 102:19]
  wire  m_21_io_x1; // @[MUL.scala 102:19]
  wire  m_21_io_x2; // @[MUL.scala 102:19]
  wire  m_21_io_x3; // @[MUL.scala 102:19]
  wire  m_21_io_s; // @[MUL.scala 102:19]
  wire  m_21_io_cout; // @[MUL.scala 102:19]
  wire  m_22_io_x1; // @[MUL.scala 102:19]
  wire  m_22_io_x2; // @[MUL.scala 102:19]
  wire  m_22_io_x3; // @[MUL.scala 102:19]
  wire  m_22_io_s; // @[MUL.scala 102:19]
  wire  m_22_io_cout; // @[MUL.scala 102:19]
  wire  m_23_io_x1; // @[MUL.scala 102:19]
  wire  m_23_io_x2; // @[MUL.scala 102:19]
  wire  m_23_io_x3; // @[MUL.scala 102:19]
  wire  m_23_io_s; // @[MUL.scala 102:19]
  wire  m_23_io_cout; // @[MUL.scala 102:19]
  wire  m_24_io_in_0; // @[MUL.scala 124:19]
  wire  m_24_io_in_1; // @[MUL.scala 124:19]
  wire  m_24_io_out_0; // @[MUL.scala 124:19]
  wire  m_24_io_out_1; // @[MUL.scala 124:19]
  wire  m_25_io_x1; // @[MUL.scala 102:19]
  wire  m_25_io_x2; // @[MUL.scala 102:19]
  wire  m_25_io_x3; // @[MUL.scala 102:19]
  wire  m_25_io_s; // @[MUL.scala 102:19]
  wire  m_25_io_cout; // @[MUL.scala 102:19]
  wire  m_26_io_in_0; // @[MUL.scala 124:19]
  wire  m_26_io_in_1; // @[MUL.scala 124:19]
  wire  m_26_io_out_0; // @[MUL.scala 124:19]
  wire  m_26_io_out_1; // @[MUL.scala 124:19]
  wire  m_27_io_x1; // @[MUL.scala 102:19]
  wire  m_27_io_x2; // @[MUL.scala 102:19]
  wire  m_27_io_x3; // @[MUL.scala 102:19]
  wire  m_27_io_s; // @[MUL.scala 102:19]
  wire  m_27_io_cout; // @[MUL.scala 102:19]
  wire  m_28_io_x1; // @[MUL.scala 102:19]
  wire  m_28_io_x2; // @[MUL.scala 102:19]
  wire  m_28_io_x3; // @[MUL.scala 102:19]
  wire  m_28_io_s; // @[MUL.scala 102:19]
  wire  m_28_io_cout; // @[MUL.scala 102:19]
  wire  m_29_io_x1; // @[MUL.scala 102:19]
  wire  m_29_io_x2; // @[MUL.scala 102:19]
  wire  m_29_io_x3; // @[MUL.scala 102:19]
  wire  m_29_io_s; // @[MUL.scala 102:19]
  wire  m_29_io_cout; // @[MUL.scala 102:19]
  wire  m_30_io_x1; // @[MUL.scala 102:19]
  wire  m_30_io_x2; // @[MUL.scala 102:19]
  wire  m_30_io_x3; // @[MUL.scala 102:19]
  wire  m_30_io_s; // @[MUL.scala 102:19]
  wire  m_30_io_cout; // @[MUL.scala 102:19]
  wire  m_31_io_x1; // @[MUL.scala 102:19]
  wire  m_31_io_x2; // @[MUL.scala 102:19]
  wire  m_31_io_x3; // @[MUL.scala 102:19]
  wire  m_31_io_s; // @[MUL.scala 102:19]
  wire  m_31_io_cout; // @[MUL.scala 102:19]
  wire  m_32_io_x1; // @[MUL.scala 102:19]
  wire  m_32_io_x2; // @[MUL.scala 102:19]
  wire  m_32_io_x3; // @[MUL.scala 102:19]
  wire  m_32_io_s; // @[MUL.scala 102:19]
  wire  m_32_io_cout; // @[MUL.scala 102:19]
  wire  m_33_io_x1; // @[MUL.scala 102:19]
  wire  m_33_io_x2; // @[MUL.scala 102:19]
  wire  m_33_io_x3; // @[MUL.scala 102:19]
  wire  m_33_io_s; // @[MUL.scala 102:19]
  wire  m_33_io_cout; // @[MUL.scala 102:19]
  wire  m_34_io_x1; // @[MUL.scala 102:19]
  wire  m_34_io_x2; // @[MUL.scala 102:19]
  wire  m_34_io_x3; // @[MUL.scala 102:19]
  wire  m_34_io_s; // @[MUL.scala 102:19]
  wire  m_34_io_cout; // @[MUL.scala 102:19]
  wire  m_35_io_x1; // @[MUL.scala 102:19]
  wire  m_35_io_x2; // @[MUL.scala 102:19]
  wire  m_35_io_x3; // @[MUL.scala 102:19]
  wire  m_35_io_s; // @[MUL.scala 102:19]
  wire  m_35_io_cout; // @[MUL.scala 102:19]
  wire  m_36_io_x1; // @[MUL.scala 102:19]
  wire  m_36_io_x2; // @[MUL.scala 102:19]
  wire  m_36_io_x3; // @[MUL.scala 102:19]
  wire  m_36_io_s; // @[MUL.scala 102:19]
  wire  m_36_io_cout; // @[MUL.scala 102:19]
  wire  m_37_io_in_0; // @[MUL.scala 124:19]
  wire  m_37_io_in_1; // @[MUL.scala 124:19]
  wire  m_37_io_out_0; // @[MUL.scala 124:19]
  wire  m_37_io_out_1; // @[MUL.scala 124:19]
  wire  m_38_io_x1; // @[MUL.scala 102:19]
  wire  m_38_io_x2; // @[MUL.scala 102:19]
  wire  m_38_io_x3; // @[MUL.scala 102:19]
  wire  m_38_io_s; // @[MUL.scala 102:19]
  wire  m_38_io_cout; // @[MUL.scala 102:19]
  wire  m_39_io_x1; // @[MUL.scala 102:19]
  wire  m_39_io_x2; // @[MUL.scala 102:19]
  wire  m_39_io_x3; // @[MUL.scala 102:19]
  wire  m_39_io_s; // @[MUL.scala 102:19]
  wire  m_39_io_cout; // @[MUL.scala 102:19]
  wire  m_40_io_in_0; // @[MUL.scala 124:19]
  wire  m_40_io_in_1; // @[MUL.scala 124:19]
  wire  m_40_io_out_0; // @[MUL.scala 124:19]
  wire  m_40_io_out_1; // @[MUL.scala 124:19]
  wire  m_41_io_x1; // @[MUL.scala 102:19]
  wire  m_41_io_x2; // @[MUL.scala 102:19]
  wire  m_41_io_x3; // @[MUL.scala 102:19]
  wire  m_41_io_s; // @[MUL.scala 102:19]
  wire  m_41_io_cout; // @[MUL.scala 102:19]
  wire  m_42_io_x1; // @[MUL.scala 102:19]
  wire  m_42_io_x2; // @[MUL.scala 102:19]
  wire  m_42_io_x3; // @[MUL.scala 102:19]
  wire  m_42_io_s; // @[MUL.scala 102:19]
  wire  m_42_io_cout; // @[MUL.scala 102:19]
  wire  m_43_io_x1; // @[MUL.scala 102:19]
  wire  m_43_io_x2; // @[MUL.scala 102:19]
  wire  m_43_io_x3; // @[MUL.scala 102:19]
  wire  m_43_io_s; // @[MUL.scala 102:19]
  wire  m_43_io_cout; // @[MUL.scala 102:19]
  wire  m_44_io_x1; // @[MUL.scala 102:19]
  wire  m_44_io_x2; // @[MUL.scala 102:19]
  wire  m_44_io_x3; // @[MUL.scala 102:19]
  wire  m_44_io_s; // @[MUL.scala 102:19]
  wire  m_44_io_cout; // @[MUL.scala 102:19]
  wire  m_45_io_x1; // @[MUL.scala 102:19]
  wire  m_45_io_x2; // @[MUL.scala 102:19]
  wire  m_45_io_x3; // @[MUL.scala 102:19]
  wire  m_45_io_s; // @[MUL.scala 102:19]
  wire  m_45_io_cout; // @[MUL.scala 102:19]
  wire  m_46_io_x1; // @[MUL.scala 102:19]
  wire  m_46_io_x2; // @[MUL.scala 102:19]
  wire  m_46_io_x3; // @[MUL.scala 102:19]
  wire  m_46_io_s; // @[MUL.scala 102:19]
  wire  m_46_io_cout; // @[MUL.scala 102:19]
  wire  m_47_io_x1; // @[MUL.scala 102:19]
  wire  m_47_io_x2; // @[MUL.scala 102:19]
  wire  m_47_io_x3; // @[MUL.scala 102:19]
  wire  m_47_io_s; // @[MUL.scala 102:19]
  wire  m_47_io_cout; // @[MUL.scala 102:19]
  wire  m_48_io_x1; // @[MUL.scala 102:19]
  wire  m_48_io_x2; // @[MUL.scala 102:19]
  wire  m_48_io_x3; // @[MUL.scala 102:19]
  wire  m_48_io_s; // @[MUL.scala 102:19]
  wire  m_48_io_cout; // @[MUL.scala 102:19]
  wire  m_49_io_x1; // @[MUL.scala 102:19]
  wire  m_49_io_x2; // @[MUL.scala 102:19]
  wire  m_49_io_x3; // @[MUL.scala 102:19]
  wire  m_49_io_s; // @[MUL.scala 102:19]
  wire  m_49_io_cout; // @[MUL.scala 102:19]
  wire  m_50_io_x1; // @[MUL.scala 102:19]
  wire  m_50_io_x2; // @[MUL.scala 102:19]
  wire  m_50_io_x3; // @[MUL.scala 102:19]
  wire  m_50_io_s; // @[MUL.scala 102:19]
  wire  m_50_io_cout; // @[MUL.scala 102:19]
  wire  m_51_io_x1; // @[MUL.scala 102:19]
  wire  m_51_io_x2; // @[MUL.scala 102:19]
  wire  m_51_io_x3; // @[MUL.scala 102:19]
  wire  m_51_io_s; // @[MUL.scala 102:19]
  wire  m_51_io_cout; // @[MUL.scala 102:19]
  wire  m_52_io_x1; // @[MUL.scala 102:19]
  wire  m_52_io_x2; // @[MUL.scala 102:19]
  wire  m_52_io_x3; // @[MUL.scala 102:19]
  wire  m_52_io_s; // @[MUL.scala 102:19]
  wire  m_52_io_cout; // @[MUL.scala 102:19]
  wire  m_53_io_x1; // @[MUL.scala 102:19]
  wire  m_53_io_x2; // @[MUL.scala 102:19]
  wire  m_53_io_x3; // @[MUL.scala 102:19]
  wire  m_53_io_s; // @[MUL.scala 102:19]
  wire  m_53_io_cout; // @[MUL.scala 102:19]
  wire  m_54_io_x1; // @[MUL.scala 102:19]
  wire  m_54_io_x2; // @[MUL.scala 102:19]
  wire  m_54_io_x3; // @[MUL.scala 102:19]
  wire  m_54_io_s; // @[MUL.scala 102:19]
  wire  m_54_io_cout; // @[MUL.scala 102:19]
  wire  m_55_io_x1; // @[MUL.scala 102:19]
  wire  m_55_io_x2; // @[MUL.scala 102:19]
  wire  m_55_io_x3; // @[MUL.scala 102:19]
  wire  m_55_io_s; // @[MUL.scala 102:19]
  wire  m_55_io_cout; // @[MUL.scala 102:19]
  wire  m_56_io_in_0; // @[MUL.scala 124:19]
  wire  m_56_io_in_1; // @[MUL.scala 124:19]
  wire  m_56_io_out_0; // @[MUL.scala 124:19]
  wire  m_56_io_out_1; // @[MUL.scala 124:19]
  wire  m_57_io_x1; // @[MUL.scala 102:19]
  wire  m_57_io_x2; // @[MUL.scala 102:19]
  wire  m_57_io_x3; // @[MUL.scala 102:19]
  wire  m_57_io_s; // @[MUL.scala 102:19]
  wire  m_57_io_cout; // @[MUL.scala 102:19]
  wire  m_58_io_x1; // @[MUL.scala 102:19]
  wire  m_58_io_x2; // @[MUL.scala 102:19]
  wire  m_58_io_x3; // @[MUL.scala 102:19]
  wire  m_58_io_s; // @[MUL.scala 102:19]
  wire  m_58_io_cout; // @[MUL.scala 102:19]
  wire  m_59_io_x1; // @[MUL.scala 102:19]
  wire  m_59_io_x2; // @[MUL.scala 102:19]
  wire  m_59_io_x3; // @[MUL.scala 102:19]
  wire  m_59_io_s; // @[MUL.scala 102:19]
  wire  m_59_io_cout; // @[MUL.scala 102:19]
  wire  m_60_io_in_0; // @[MUL.scala 124:19]
  wire  m_60_io_in_1; // @[MUL.scala 124:19]
  wire  m_60_io_out_0; // @[MUL.scala 124:19]
  wire  m_60_io_out_1; // @[MUL.scala 124:19]
  wire  m_61_io_x1; // @[MUL.scala 102:19]
  wire  m_61_io_x2; // @[MUL.scala 102:19]
  wire  m_61_io_x3; // @[MUL.scala 102:19]
  wire  m_61_io_s; // @[MUL.scala 102:19]
  wire  m_61_io_cout; // @[MUL.scala 102:19]
  wire  m_62_io_x1; // @[MUL.scala 102:19]
  wire  m_62_io_x2; // @[MUL.scala 102:19]
  wire  m_62_io_x3; // @[MUL.scala 102:19]
  wire  m_62_io_s; // @[MUL.scala 102:19]
  wire  m_62_io_cout; // @[MUL.scala 102:19]
  wire  m_63_io_x1; // @[MUL.scala 102:19]
  wire  m_63_io_x2; // @[MUL.scala 102:19]
  wire  m_63_io_x3; // @[MUL.scala 102:19]
  wire  m_63_io_s; // @[MUL.scala 102:19]
  wire  m_63_io_cout; // @[MUL.scala 102:19]
  wire  m_64_io_x1; // @[MUL.scala 102:19]
  wire  m_64_io_x2; // @[MUL.scala 102:19]
  wire  m_64_io_x3; // @[MUL.scala 102:19]
  wire  m_64_io_s; // @[MUL.scala 102:19]
  wire  m_64_io_cout; // @[MUL.scala 102:19]
  wire  m_65_io_x1; // @[MUL.scala 102:19]
  wire  m_65_io_x2; // @[MUL.scala 102:19]
  wire  m_65_io_x3; // @[MUL.scala 102:19]
  wire  m_65_io_s; // @[MUL.scala 102:19]
  wire  m_65_io_cout; // @[MUL.scala 102:19]
  wire  m_66_io_x1; // @[MUL.scala 102:19]
  wire  m_66_io_x2; // @[MUL.scala 102:19]
  wire  m_66_io_x3; // @[MUL.scala 102:19]
  wire  m_66_io_s; // @[MUL.scala 102:19]
  wire  m_66_io_cout; // @[MUL.scala 102:19]
  wire  m_67_io_x1; // @[MUL.scala 102:19]
  wire  m_67_io_x2; // @[MUL.scala 102:19]
  wire  m_67_io_x3; // @[MUL.scala 102:19]
  wire  m_67_io_s; // @[MUL.scala 102:19]
  wire  m_67_io_cout; // @[MUL.scala 102:19]
  wire  m_68_io_x1; // @[MUL.scala 102:19]
  wire  m_68_io_x2; // @[MUL.scala 102:19]
  wire  m_68_io_x3; // @[MUL.scala 102:19]
  wire  m_68_io_s; // @[MUL.scala 102:19]
  wire  m_68_io_cout; // @[MUL.scala 102:19]
  wire  m_69_io_x1; // @[MUL.scala 102:19]
  wire  m_69_io_x2; // @[MUL.scala 102:19]
  wire  m_69_io_x3; // @[MUL.scala 102:19]
  wire  m_69_io_s; // @[MUL.scala 102:19]
  wire  m_69_io_cout; // @[MUL.scala 102:19]
  wire  m_70_io_x1; // @[MUL.scala 102:19]
  wire  m_70_io_x2; // @[MUL.scala 102:19]
  wire  m_70_io_x3; // @[MUL.scala 102:19]
  wire  m_70_io_s; // @[MUL.scala 102:19]
  wire  m_70_io_cout; // @[MUL.scala 102:19]
  wire  m_71_io_x1; // @[MUL.scala 102:19]
  wire  m_71_io_x2; // @[MUL.scala 102:19]
  wire  m_71_io_x3; // @[MUL.scala 102:19]
  wire  m_71_io_s; // @[MUL.scala 102:19]
  wire  m_71_io_cout; // @[MUL.scala 102:19]
  wire  m_72_io_x1; // @[MUL.scala 102:19]
  wire  m_72_io_x2; // @[MUL.scala 102:19]
  wire  m_72_io_x3; // @[MUL.scala 102:19]
  wire  m_72_io_s; // @[MUL.scala 102:19]
  wire  m_72_io_cout; // @[MUL.scala 102:19]
  wire  m_73_io_x1; // @[MUL.scala 102:19]
  wire  m_73_io_x2; // @[MUL.scala 102:19]
  wire  m_73_io_x3; // @[MUL.scala 102:19]
  wire  m_73_io_s; // @[MUL.scala 102:19]
  wire  m_73_io_cout; // @[MUL.scala 102:19]
  wire  m_74_io_x1; // @[MUL.scala 102:19]
  wire  m_74_io_x2; // @[MUL.scala 102:19]
  wire  m_74_io_x3; // @[MUL.scala 102:19]
  wire  m_74_io_s; // @[MUL.scala 102:19]
  wire  m_74_io_cout; // @[MUL.scala 102:19]
  wire  m_75_io_x1; // @[MUL.scala 102:19]
  wire  m_75_io_x2; // @[MUL.scala 102:19]
  wire  m_75_io_x3; // @[MUL.scala 102:19]
  wire  m_75_io_s; // @[MUL.scala 102:19]
  wire  m_75_io_cout; // @[MUL.scala 102:19]
  wire  m_76_io_x1; // @[MUL.scala 102:19]
  wire  m_76_io_x2; // @[MUL.scala 102:19]
  wire  m_76_io_x3; // @[MUL.scala 102:19]
  wire  m_76_io_s; // @[MUL.scala 102:19]
  wire  m_76_io_cout; // @[MUL.scala 102:19]
  wire  m_77_io_x1; // @[MUL.scala 102:19]
  wire  m_77_io_x2; // @[MUL.scala 102:19]
  wire  m_77_io_x3; // @[MUL.scala 102:19]
  wire  m_77_io_s; // @[MUL.scala 102:19]
  wire  m_77_io_cout; // @[MUL.scala 102:19]
  wire  m_78_io_x1; // @[MUL.scala 102:19]
  wire  m_78_io_x2; // @[MUL.scala 102:19]
  wire  m_78_io_x3; // @[MUL.scala 102:19]
  wire  m_78_io_s; // @[MUL.scala 102:19]
  wire  m_78_io_cout; // @[MUL.scala 102:19]
  wire  m_79_io_x1; // @[MUL.scala 102:19]
  wire  m_79_io_x2; // @[MUL.scala 102:19]
  wire  m_79_io_x3; // @[MUL.scala 102:19]
  wire  m_79_io_s; // @[MUL.scala 102:19]
  wire  m_79_io_cout; // @[MUL.scala 102:19]
  wire  m_80_io_x1; // @[MUL.scala 102:19]
  wire  m_80_io_x2; // @[MUL.scala 102:19]
  wire  m_80_io_x3; // @[MUL.scala 102:19]
  wire  m_80_io_s; // @[MUL.scala 102:19]
  wire  m_80_io_cout; // @[MUL.scala 102:19]
  wire  m_81_io_in_0; // @[MUL.scala 124:19]
  wire  m_81_io_in_1; // @[MUL.scala 124:19]
  wire  m_81_io_out_0; // @[MUL.scala 124:19]
  wire  m_81_io_out_1; // @[MUL.scala 124:19]
  wire  m_82_io_x1; // @[MUL.scala 102:19]
  wire  m_82_io_x2; // @[MUL.scala 102:19]
  wire  m_82_io_x3; // @[MUL.scala 102:19]
  wire  m_82_io_s; // @[MUL.scala 102:19]
  wire  m_82_io_cout; // @[MUL.scala 102:19]
  wire  m_83_io_x1; // @[MUL.scala 102:19]
  wire  m_83_io_x2; // @[MUL.scala 102:19]
  wire  m_83_io_x3; // @[MUL.scala 102:19]
  wire  m_83_io_s; // @[MUL.scala 102:19]
  wire  m_83_io_cout; // @[MUL.scala 102:19]
  wire  m_84_io_x1; // @[MUL.scala 102:19]
  wire  m_84_io_x2; // @[MUL.scala 102:19]
  wire  m_84_io_x3; // @[MUL.scala 102:19]
  wire  m_84_io_s; // @[MUL.scala 102:19]
  wire  m_84_io_cout; // @[MUL.scala 102:19]
  wire  m_85_io_x1; // @[MUL.scala 102:19]
  wire  m_85_io_x2; // @[MUL.scala 102:19]
  wire  m_85_io_x3; // @[MUL.scala 102:19]
  wire  m_85_io_s; // @[MUL.scala 102:19]
  wire  m_85_io_cout; // @[MUL.scala 102:19]
  wire  m_86_io_in_0; // @[MUL.scala 124:19]
  wire  m_86_io_in_1; // @[MUL.scala 124:19]
  wire  m_86_io_out_0; // @[MUL.scala 124:19]
  wire  m_86_io_out_1; // @[MUL.scala 124:19]
  wire  m_87_io_x1; // @[MUL.scala 102:19]
  wire  m_87_io_x2; // @[MUL.scala 102:19]
  wire  m_87_io_x3; // @[MUL.scala 102:19]
  wire  m_87_io_s; // @[MUL.scala 102:19]
  wire  m_87_io_cout; // @[MUL.scala 102:19]
  wire  m_88_io_x1; // @[MUL.scala 102:19]
  wire  m_88_io_x2; // @[MUL.scala 102:19]
  wire  m_88_io_x3; // @[MUL.scala 102:19]
  wire  m_88_io_s; // @[MUL.scala 102:19]
  wire  m_88_io_cout; // @[MUL.scala 102:19]
  wire  m_89_io_x1; // @[MUL.scala 102:19]
  wire  m_89_io_x2; // @[MUL.scala 102:19]
  wire  m_89_io_x3; // @[MUL.scala 102:19]
  wire  m_89_io_s; // @[MUL.scala 102:19]
  wire  m_89_io_cout; // @[MUL.scala 102:19]
  wire  m_90_io_x1; // @[MUL.scala 102:19]
  wire  m_90_io_x2; // @[MUL.scala 102:19]
  wire  m_90_io_x3; // @[MUL.scala 102:19]
  wire  m_90_io_s; // @[MUL.scala 102:19]
  wire  m_90_io_cout; // @[MUL.scala 102:19]
  wire  m_91_io_x1; // @[MUL.scala 102:19]
  wire  m_91_io_x2; // @[MUL.scala 102:19]
  wire  m_91_io_x3; // @[MUL.scala 102:19]
  wire  m_91_io_s; // @[MUL.scala 102:19]
  wire  m_91_io_cout; // @[MUL.scala 102:19]
  wire  m_92_io_x1; // @[MUL.scala 102:19]
  wire  m_92_io_x2; // @[MUL.scala 102:19]
  wire  m_92_io_x3; // @[MUL.scala 102:19]
  wire  m_92_io_s; // @[MUL.scala 102:19]
  wire  m_92_io_cout; // @[MUL.scala 102:19]
  wire  m_93_io_x1; // @[MUL.scala 102:19]
  wire  m_93_io_x2; // @[MUL.scala 102:19]
  wire  m_93_io_x3; // @[MUL.scala 102:19]
  wire  m_93_io_s; // @[MUL.scala 102:19]
  wire  m_93_io_cout; // @[MUL.scala 102:19]
  wire  m_94_io_x1; // @[MUL.scala 102:19]
  wire  m_94_io_x2; // @[MUL.scala 102:19]
  wire  m_94_io_x3; // @[MUL.scala 102:19]
  wire  m_94_io_s; // @[MUL.scala 102:19]
  wire  m_94_io_cout; // @[MUL.scala 102:19]
  wire  m_95_io_x1; // @[MUL.scala 102:19]
  wire  m_95_io_x2; // @[MUL.scala 102:19]
  wire  m_95_io_x3; // @[MUL.scala 102:19]
  wire  m_95_io_s; // @[MUL.scala 102:19]
  wire  m_95_io_cout; // @[MUL.scala 102:19]
  wire  m_96_io_x1; // @[MUL.scala 102:19]
  wire  m_96_io_x2; // @[MUL.scala 102:19]
  wire  m_96_io_x3; // @[MUL.scala 102:19]
  wire  m_96_io_s; // @[MUL.scala 102:19]
  wire  m_96_io_cout; // @[MUL.scala 102:19]
  wire  m_97_io_x1; // @[MUL.scala 102:19]
  wire  m_97_io_x2; // @[MUL.scala 102:19]
  wire  m_97_io_x3; // @[MUL.scala 102:19]
  wire  m_97_io_s; // @[MUL.scala 102:19]
  wire  m_97_io_cout; // @[MUL.scala 102:19]
  wire  m_98_io_x1; // @[MUL.scala 102:19]
  wire  m_98_io_x2; // @[MUL.scala 102:19]
  wire  m_98_io_x3; // @[MUL.scala 102:19]
  wire  m_98_io_s; // @[MUL.scala 102:19]
  wire  m_98_io_cout; // @[MUL.scala 102:19]
  wire  m_99_io_x1; // @[MUL.scala 102:19]
  wire  m_99_io_x2; // @[MUL.scala 102:19]
  wire  m_99_io_x3; // @[MUL.scala 102:19]
  wire  m_99_io_s; // @[MUL.scala 102:19]
  wire  m_99_io_cout; // @[MUL.scala 102:19]
  wire  m_100_io_x1; // @[MUL.scala 102:19]
  wire  m_100_io_x2; // @[MUL.scala 102:19]
  wire  m_100_io_x3; // @[MUL.scala 102:19]
  wire  m_100_io_s; // @[MUL.scala 102:19]
  wire  m_100_io_cout; // @[MUL.scala 102:19]
  wire  m_101_io_x1; // @[MUL.scala 102:19]
  wire  m_101_io_x2; // @[MUL.scala 102:19]
  wire  m_101_io_x3; // @[MUL.scala 102:19]
  wire  m_101_io_s; // @[MUL.scala 102:19]
  wire  m_101_io_cout; // @[MUL.scala 102:19]
  wire  m_102_io_x1; // @[MUL.scala 102:19]
  wire  m_102_io_x2; // @[MUL.scala 102:19]
  wire  m_102_io_x3; // @[MUL.scala 102:19]
  wire  m_102_io_s; // @[MUL.scala 102:19]
  wire  m_102_io_cout; // @[MUL.scala 102:19]
  wire  m_103_io_x1; // @[MUL.scala 102:19]
  wire  m_103_io_x2; // @[MUL.scala 102:19]
  wire  m_103_io_x3; // @[MUL.scala 102:19]
  wire  m_103_io_s; // @[MUL.scala 102:19]
  wire  m_103_io_cout; // @[MUL.scala 102:19]
  wire  m_104_io_x1; // @[MUL.scala 102:19]
  wire  m_104_io_x2; // @[MUL.scala 102:19]
  wire  m_104_io_x3; // @[MUL.scala 102:19]
  wire  m_104_io_s; // @[MUL.scala 102:19]
  wire  m_104_io_cout; // @[MUL.scala 102:19]
  wire  m_105_io_x1; // @[MUL.scala 102:19]
  wire  m_105_io_x2; // @[MUL.scala 102:19]
  wire  m_105_io_x3; // @[MUL.scala 102:19]
  wire  m_105_io_s; // @[MUL.scala 102:19]
  wire  m_105_io_cout; // @[MUL.scala 102:19]
  wire  m_106_io_x1; // @[MUL.scala 102:19]
  wire  m_106_io_x2; // @[MUL.scala 102:19]
  wire  m_106_io_x3; // @[MUL.scala 102:19]
  wire  m_106_io_s; // @[MUL.scala 102:19]
  wire  m_106_io_cout; // @[MUL.scala 102:19]
  wire  m_107_io_x1; // @[MUL.scala 102:19]
  wire  m_107_io_x2; // @[MUL.scala 102:19]
  wire  m_107_io_x3; // @[MUL.scala 102:19]
  wire  m_107_io_s; // @[MUL.scala 102:19]
  wire  m_107_io_cout; // @[MUL.scala 102:19]
  wire  m_108_io_x1; // @[MUL.scala 102:19]
  wire  m_108_io_x2; // @[MUL.scala 102:19]
  wire  m_108_io_x3; // @[MUL.scala 102:19]
  wire  m_108_io_s; // @[MUL.scala 102:19]
  wire  m_108_io_cout; // @[MUL.scala 102:19]
  wire  m_109_io_x1; // @[MUL.scala 102:19]
  wire  m_109_io_x2; // @[MUL.scala 102:19]
  wire  m_109_io_x3; // @[MUL.scala 102:19]
  wire  m_109_io_s; // @[MUL.scala 102:19]
  wire  m_109_io_cout; // @[MUL.scala 102:19]
  wire  m_110_io_x1; // @[MUL.scala 102:19]
  wire  m_110_io_x2; // @[MUL.scala 102:19]
  wire  m_110_io_x3; // @[MUL.scala 102:19]
  wire  m_110_io_s; // @[MUL.scala 102:19]
  wire  m_110_io_cout; // @[MUL.scala 102:19]
  wire  m_111_io_x1; // @[MUL.scala 102:19]
  wire  m_111_io_x2; // @[MUL.scala 102:19]
  wire  m_111_io_x3; // @[MUL.scala 102:19]
  wire  m_111_io_s; // @[MUL.scala 102:19]
  wire  m_111_io_cout; // @[MUL.scala 102:19]
  wire  m_112_io_in_0; // @[MUL.scala 124:19]
  wire  m_112_io_in_1; // @[MUL.scala 124:19]
  wire  m_112_io_out_0; // @[MUL.scala 124:19]
  wire  m_112_io_out_1; // @[MUL.scala 124:19]
  wire  m_113_io_x1; // @[MUL.scala 102:19]
  wire  m_113_io_x2; // @[MUL.scala 102:19]
  wire  m_113_io_x3; // @[MUL.scala 102:19]
  wire  m_113_io_s; // @[MUL.scala 102:19]
  wire  m_113_io_cout; // @[MUL.scala 102:19]
  wire  m_114_io_x1; // @[MUL.scala 102:19]
  wire  m_114_io_x2; // @[MUL.scala 102:19]
  wire  m_114_io_x3; // @[MUL.scala 102:19]
  wire  m_114_io_s; // @[MUL.scala 102:19]
  wire  m_114_io_cout; // @[MUL.scala 102:19]
  wire  m_115_io_x1; // @[MUL.scala 102:19]
  wire  m_115_io_x2; // @[MUL.scala 102:19]
  wire  m_115_io_x3; // @[MUL.scala 102:19]
  wire  m_115_io_s; // @[MUL.scala 102:19]
  wire  m_115_io_cout; // @[MUL.scala 102:19]
  wire  m_116_io_x1; // @[MUL.scala 102:19]
  wire  m_116_io_x2; // @[MUL.scala 102:19]
  wire  m_116_io_x3; // @[MUL.scala 102:19]
  wire  m_116_io_s; // @[MUL.scala 102:19]
  wire  m_116_io_cout; // @[MUL.scala 102:19]
  wire  m_117_io_x1; // @[MUL.scala 102:19]
  wire  m_117_io_x2; // @[MUL.scala 102:19]
  wire  m_117_io_x3; // @[MUL.scala 102:19]
  wire  m_117_io_s; // @[MUL.scala 102:19]
  wire  m_117_io_cout; // @[MUL.scala 102:19]
  wire  m_118_io_in_0; // @[MUL.scala 124:19]
  wire  m_118_io_in_1; // @[MUL.scala 124:19]
  wire  m_118_io_out_0; // @[MUL.scala 124:19]
  wire  m_118_io_out_1; // @[MUL.scala 124:19]
  wire  m_119_io_x1; // @[MUL.scala 102:19]
  wire  m_119_io_x2; // @[MUL.scala 102:19]
  wire  m_119_io_x3; // @[MUL.scala 102:19]
  wire  m_119_io_s; // @[MUL.scala 102:19]
  wire  m_119_io_cout; // @[MUL.scala 102:19]
  wire  m_120_io_x1; // @[MUL.scala 102:19]
  wire  m_120_io_x2; // @[MUL.scala 102:19]
  wire  m_120_io_x3; // @[MUL.scala 102:19]
  wire  m_120_io_s; // @[MUL.scala 102:19]
  wire  m_120_io_cout; // @[MUL.scala 102:19]
  wire  m_121_io_x1; // @[MUL.scala 102:19]
  wire  m_121_io_x2; // @[MUL.scala 102:19]
  wire  m_121_io_x3; // @[MUL.scala 102:19]
  wire  m_121_io_s; // @[MUL.scala 102:19]
  wire  m_121_io_cout; // @[MUL.scala 102:19]
  wire  m_122_io_x1; // @[MUL.scala 102:19]
  wire  m_122_io_x2; // @[MUL.scala 102:19]
  wire  m_122_io_x3; // @[MUL.scala 102:19]
  wire  m_122_io_s; // @[MUL.scala 102:19]
  wire  m_122_io_cout; // @[MUL.scala 102:19]
  wire  m_123_io_x1; // @[MUL.scala 102:19]
  wire  m_123_io_x2; // @[MUL.scala 102:19]
  wire  m_123_io_x3; // @[MUL.scala 102:19]
  wire  m_123_io_s; // @[MUL.scala 102:19]
  wire  m_123_io_cout; // @[MUL.scala 102:19]
  wire  m_124_io_in_0; // @[MUL.scala 124:19]
  wire  m_124_io_in_1; // @[MUL.scala 124:19]
  wire  m_124_io_out_0; // @[MUL.scala 124:19]
  wire  m_124_io_out_1; // @[MUL.scala 124:19]
  wire  m_125_io_x1; // @[MUL.scala 102:19]
  wire  m_125_io_x2; // @[MUL.scala 102:19]
  wire  m_125_io_x3; // @[MUL.scala 102:19]
  wire  m_125_io_s; // @[MUL.scala 102:19]
  wire  m_125_io_cout; // @[MUL.scala 102:19]
  wire  m_126_io_x1; // @[MUL.scala 102:19]
  wire  m_126_io_x2; // @[MUL.scala 102:19]
  wire  m_126_io_x3; // @[MUL.scala 102:19]
  wire  m_126_io_s; // @[MUL.scala 102:19]
  wire  m_126_io_cout; // @[MUL.scala 102:19]
  wire  m_127_io_x1; // @[MUL.scala 102:19]
  wire  m_127_io_x2; // @[MUL.scala 102:19]
  wire  m_127_io_x3; // @[MUL.scala 102:19]
  wire  m_127_io_s; // @[MUL.scala 102:19]
  wire  m_127_io_cout; // @[MUL.scala 102:19]
  wire  m_128_io_x1; // @[MUL.scala 102:19]
  wire  m_128_io_x2; // @[MUL.scala 102:19]
  wire  m_128_io_x3; // @[MUL.scala 102:19]
  wire  m_128_io_s; // @[MUL.scala 102:19]
  wire  m_128_io_cout; // @[MUL.scala 102:19]
  wire  m_129_io_x1; // @[MUL.scala 102:19]
  wire  m_129_io_x2; // @[MUL.scala 102:19]
  wire  m_129_io_x3; // @[MUL.scala 102:19]
  wire  m_129_io_s; // @[MUL.scala 102:19]
  wire  m_129_io_cout; // @[MUL.scala 102:19]
  wire  m_130_io_in_0; // @[MUL.scala 124:19]
  wire  m_130_io_in_1; // @[MUL.scala 124:19]
  wire  m_130_io_out_0; // @[MUL.scala 124:19]
  wire  m_130_io_out_1; // @[MUL.scala 124:19]
  wire  m_131_io_x1; // @[MUL.scala 102:19]
  wire  m_131_io_x2; // @[MUL.scala 102:19]
  wire  m_131_io_x3; // @[MUL.scala 102:19]
  wire  m_131_io_s; // @[MUL.scala 102:19]
  wire  m_131_io_cout; // @[MUL.scala 102:19]
  wire  m_132_io_x1; // @[MUL.scala 102:19]
  wire  m_132_io_x2; // @[MUL.scala 102:19]
  wire  m_132_io_x3; // @[MUL.scala 102:19]
  wire  m_132_io_s; // @[MUL.scala 102:19]
  wire  m_132_io_cout; // @[MUL.scala 102:19]
  wire  m_133_io_x1; // @[MUL.scala 102:19]
  wire  m_133_io_x2; // @[MUL.scala 102:19]
  wire  m_133_io_x3; // @[MUL.scala 102:19]
  wire  m_133_io_s; // @[MUL.scala 102:19]
  wire  m_133_io_cout; // @[MUL.scala 102:19]
  wire  m_134_io_x1; // @[MUL.scala 102:19]
  wire  m_134_io_x2; // @[MUL.scala 102:19]
  wire  m_134_io_x3; // @[MUL.scala 102:19]
  wire  m_134_io_s; // @[MUL.scala 102:19]
  wire  m_134_io_cout; // @[MUL.scala 102:19]
  wire  m_135_io_x1; // @[MUL.scala 102:19]
  wire  m_135_io_x2; // @[MUL.scala 102:19]
  wire  m_135_io_x3; // @[MUL.scala 102:19]
  wire  m_135_io_s; // @[MUL.scala 102:19]
  wire  m_135_io_cout; // @[MUL.scala 102:19]
  wire  m_136_io_in_0; // @[MUL.scala 124:19]
  wire  m_136_io_in_1; // @[MUL.scala 124:19]
  wire  m_136_io_out_0; // @[MUL.scala 124:19]
  wire  m_136_io_out_1; // @[MUL.scala 124:19]
  wire  m_137_io_x1; // @[MUL.scala 102:19]
  wire  m_137_io_x2; // @[MUL.scala 102:19]
  wire  m_137_io_x3; // @[MUL.scala 102:19]
  wire  m_137_io_s; // @[MUL.scala 102:19]
  wire  m_137_io_cout; // @[MUL.scala 102:19]
  wire  m_138_io_x1; // @[MUL.scala 102:19]
  wire  m_138_io_x2; // @[MUL.scala 102:19]
  wire  m_138_io_x3; // @[MUL.scala 102:19]
  wire  m_138_io_s; // @[MUL.scala 102:19]
  wire  m_138_io_cout; // @[MUL.scala 102:19]
  wire  m_139_io_x1; // @[MUL.scala 102:19]
  wire  m_139_io_x2; // @[MUL.scala 102:19]
  wire  m_139_io_x3; // @[MUL.scala 102:19]
  wire  m_139_io_s; // @[MUL.scala 102:19]
  wire  m_139_io_cout; // @[MUL.scala 102:19]
  wire  m_140_io_x1; // @[MUL.scala 102:19]
  wire  m_140_io_x2; // @[MUL.scala 102:19]
  wire  m_140_io_x3; // @[MUL.scala 102:19]
  wire  m_140_io_s; // @[MUL.scala 102:19]
  wire  m_140_io_cout; // @[MUL.scala 102:19]
  wire  m_141_io_x1; // @[MUL.scala 102:19]
  wire  m_141_io_x2; // @[MUL.scala 102:19]
  wire  m_141_io_x3; // @[MUL.scala 102:19]
  wire  m_141_io_s; // @[MUL.scala 102:19]
  wire  m_141_io_cout; // @[MUL.scala 102:19]
  wire  m_142_io_in_0; // @[MUL.scala 124:19]
  wire  m_142_io_in_1; // @[MUL.scala 124:19]
  wire  m_142_io_out_0; // @[MUL.scala 124:19]
  wire  m_142_io_out_1; // @[MUL.scala 124:19]
  wire  m_143_io_x1; // @[MUL.scala 102:19]
  wire  m_143_io_x2; // @[MUL.scala 102:19]
  wire  m_143_io_x3; // @[MUL.scala 102:19]
  wire  m_143_io_s; // @[MUL.scala 102:19]
  wire  m_143_io_cout; // @[MUL.scala 102:19]
  wire  m_144_io_x1; // @[MUL.scala 102:19]
  wire  m_144_io_x2; // @[MUL.scala 102:19]
  wire  m_144_io_x3; // @[MUL.scala 102:19]
  wire  m_144_io_s; // @[MUL.scala 102:19]
  wire  m_144_io_cout; // @[MUL.scala 102:19]
  wire  m_145_io_x1; // @[MUL.scala 102:19]
  wire  m_145_io_x2; // @[MUL.scala 102:19]
  wire  m_145_io_x3; // @[MUL.scala 102:19]
  wire  m_145_io_s; // @[MUL.scala 102:19]
  wire  m_145_io_cout; // @[MUL.scala 102:19]
  wire  m_146_io_x1; // @[MUL.scala 102:19]
  wire  m_146_io_x2; // @[MUL.scala 102:19]
  wire  m_146_io_x3; // @[MUL.scala 102:19]
  wire  m_146_io_s; // @[MUL.scala 102:19]
  wire  m_146_io_cout; // @[MUL.scala 102:19]
  wire  m_147_io_x1; // @[MUL.scala 102:19]
  wire  m_147_io_x2; // @[MUL.scala 102:19]
  wire  m_147_io_x3; // @[MUL.scala 102:19]
  wire  m_147_io_s; // @[MUL.scala 102:19]
  wire  m_147_io_cout; // @[MUL.scala 102:19]
  wire  m_148_io_in_0; // @[MUL.scala 124:19]
  wire  m_148_io_in_1; // @[MUL.scala 124:19]
  wire  m_148_io_out_0; // @[MUL.scala 124:19]
  wire  m_148_io_out_1; // @[MUL.scala 124:19]
  wire  m_149_io_x1; // @[MUL.scala 102:19]
  wire  m_149_io_x2; // @[MUL.scala 102:19]
  wire  m_149_io_x3; // @[MUL.scala 102:19]
  wire  m_149_io_s; // @[MUL.scala 102:19]
  wire  m_149_io_cout; // @[MUL.scala 102:19]
  wire  m_150_io_x1; // @[MUL.scala 102:19]
  wire  m_150_io_x2; // @[MUL.scala 102:19]
  wire  m_150_io_x3; // @[MUL.scala 102:19]
  wire  m_150_io_s; // @[MUL.scala 102:19]
  wire  m_150_io_cout; // @[MUL.scala 102:19]
  wire  m_151_io_x1; // @[MUL.scala 102:19]
  wire  m_151_io_x2; // @[MUL.scala 102:19]
  wire  m_151_io_x3; // @[MUL.scala 102:19]
  wire  m_151_io_s; // @[MUL.scala 102:19]
  wire  m_151_io_cout; // @[MUL.scala 102:19]
  wire  m_152_io_x1; // @[MUL.scala 102:19]
  wire  m_152_io_x2; // @[MUL.scala 102:19]
  wire  m_152_io_x3; // @[MUL.scala 102:19]
  wire  m_152_io_s; // @[MUL.scala 102:19]
  wire  m_152_io_cout; // @[MUL.scala 102:19]
  wire  m_153_io_x1; // @[MUL.scala 102:19]
  wire  m_153_io_x2; // @[MUL.scala 102:19]
  wire  m_153_io_x3; // @[MUL.scala 102:19]
  wire  m_153_io_s; // @[MUL.scala 102:19]
  wire  m_153_io_cout; // @[MUL.scala 102:19]
  wire  m_154_io_x1; // @[MUL.scala 102:19]
  wire  m_154_io_x2; // @[MUL.scala 102:19]
  wire  m_154_io_x3; // @[MUL.scala 102:19]
  wire  m_154_io_s; // @[MUL.scala 102:19]
  wire  m_154_io_cout; // @[MUL.scala 102:19]
  wire  m_155_io_x1; // @[MUL.scala 102:19]
  wire  m_155_io_x2; // @[MUL.scala 102:19]
  wire  m_155_io_x3; // @[MUL.scala 102:19]
  wire  m_155_io_s; // @[MUL.scala 102:19]
  wire  m_155_io_cout; // @[MUL.scala 102:19]
  wire  m_156_io_x1; // @[MUL.scala 102:19]
  wire  m_156_io_x2; // @[MUL.scala 102:19]
  wire  m_156_io_x3; // @[MUL.scala 102:19]
  wire  m_156_io_s; // @[MUL.scala 102:19]
  wire  m_156_io_cout; // @[MUL.scala 102:19]
  wire  m_157_io_x1; // @[MUL.scala 102:19]
  wire  m_157_io_x2; // @[MUL.scala 102:19]
  wire  m_157_io_x3; // @[MUL.scala 102:19]
  wire  m_157_io_s; // @[MUL.scala 102:19]
  wire  m_157_io_cout; // @[MUL.scala 102:19]
  wire  m_158_io_x1; // @[MUL.scala 102:19]
  wire  m_158_io_x2; // @[MUL.scala 102:19]
  wire  m_158_io_x3; // @[MUL.scala 102:19]
  wire  m_158_io_s; // @[MUL.scala 102:19]
  wire  m_158_io_cout; // @[MUL.scala 102:19]
  wire  m_159_io_x1; // @[MUL.scala 102:19]
  wire  m_159_io_x2; // @[MUL.scala 102:19]
  wire  m_159_io_x3; // @[MUL.scala 102:19]
  wire  m_159_io_s; // @[MUL.scala 102:19]
  wire  m_159_io_cout; // @[MUL.scala 102:19]
  wire  m_160_io_x1; // @[MUL.scala 102:19]
  wire  m_160_io_x2; // @[MUL.scala 102:19]
  wire  m_160_io_x3; // @[MUL.scala 102:19]
  wire  m_160_io_s; // @[MUL.scala 102:19]
  wire  m_160_io_cout; // @[MUL.scala 102:19]
  wire  m_161_io_x1; // @[MUL.scala 102:19]
  wire  m_161_io_x2; // @[MUL.scala 102:19]
  wire  m_161_io_x3; // @[MUL.scala 102:19]
  wire  m_161_io_s; // @[MUL.scala 102:19]
  wire  m_161_io_cout; // @[MUL.scala 102:19]
  wire  m_162_io_x1; // @[MUL.scala 102:19]
  wire  m_162_io_x2; // @[MUL.scala 102:19]
  wire  m_162_io_x3; // @[MUL.scala 102:19]
  wire  m_162_io_s; // @[MUL.scala 102:19]
  wire  m_162_io_cout; // @[MUL.scala 102:19]
  wire  m_163_io_x1; // @[MUL.scala 102:19]
  wire  m_163_io_x2; // @[MUL.scala 102:19]
  wire  m_163_io_x3; // @[MUL.scala 102:19]
  wire  m_163_io_s; // @[MUL.scala 102:19]
  wire  m_163_io_cout; // @[MUL.scala 102:19]
  wire  m_164_io_x1; // @[MUL.scala 102:19]
  wire  m_164_io_x2; // @[MUL.scala 102:19]
  wire  m_164_io_x3; // @[MUL.scala 102:19]
  wire  m_164_io_s; // @[MUL.scala 102:19]
  wire  m_164_io_cout; // @[MUL.scala 102:19]
  wire  m_165_io_x1; // @[MUL.scala 102:19]
  wire  m_165_io_x2; // @[MUL.scala 102:19]
  wire  m_165_io_x3; // @[MUL.scala 102:19]
  wire  m_165_io_s; // @[MUL.scala 102:19]
  wire  m_165_io_cout; // @[MUL.scala 102:19]
  wire  m_166_io_x1; // @[MUL.scala 102:19]
  wire  m_166_io_x2; // @[MUL.scala 102:19]
  wire  m_166_io_x3; // @[MUL.scala 102:19]
  wire  m_166_io_s; // @[MUL.scala 102:19]
  wire  m_166_io_cout; // @[MUL.scala 102:19]
  wire  m_167_io_x1; // @[MUL.scala 102:19]
  wire  m_167_io_x2; // @[MUL.scala 102:19]
  wire  m_167_io_x3; // @[MUL.scala 102:19]
  wire  m_167_io_s; // @[MUL.scala 102:19]
  wire  m_167_io_cout; // @[MUL.scala 102:19]
  wire  m_168_io_in_0; // @[MUL.scala 124:19]
  wire  m_168_io_in_1; // @[MUL.scala 124:19]
  wire  m_168_io_out_0; // @[MUL.scala 124:19]
  wire  m_168_io_out_1; // @[MUL.scala 124:19]
  wire  m_169_io_x1; // @[MUL.scala 102:19]
  wire  m_169_io_x2; // @[MUL.scala 102:19]
  wire  m_169_io_x3; // @[MUL.scala 102:19]
  wire  m_169_io_s; // @[MUL.scala 102:19]
  wire  m_169_io_cout; // @[MUL.scala 102:19]
  wire  m_170_io_x1; // @[MUL.scala 102:19]
  wire  m_170_io_x2; // @[MUL.scala 102:19]
  wire  m_170_io_x3; // @[MUL.scala 102:19]
  wire  m_170_io_s; // @[MUL.scala 102:19]
  wire  m_170_io_cout; // @[MUL.scala 102:19]
  wire  m_171_io_x1; // @[MUL.scala 102:19]
  wire  m_171_io_x2; // @[MUL.scala 102:19]
  wire  m_171_io_x3; // @[MUL.scala 102:19]
  wire  m_171_io_s; // @[MUL.scala 102:19]
  wire  m_171_io_cout; // @[MUL.scala 102:19]
  wire  m_172_io_x1; // @[MUL.scala 102:19]
  wire  m_172_io_x2; // @[MUL.scala 102:19]
  wire  m_172_io_x3; // @[MUL.scala 102:19]
  wire  m_172_io_s; // @[MUL.scala 102:19]
  wire  m_172_io_cout; // @[MUL.scala 102:19]
  wire  m_173_io_in_0; // @[MUL.scala 124:19]
  wire  m_173_io_in_1; // @[MUL.scala 124:19]
  wire  m_173_io_out_0; // @[MUL.scala 124:19]
  wire  m_173_io_out_1; // @[MUL.scala 124:19]
  wire  m_174_io_x1; // @[MUL.scala 102:19]
  wire  m_174_io_x2; // @[MUL.scala 102:19]
  wire  m_174_io_x3; // @[MUL.scala 102:19]
  wire  m_174_io_s; // @[MUL.scala 102:19]
  wire  m_174_io_cout; // @[MUL.scala 102:19]
  wire  m_175_io_x1; // @[MUL.scala 102:19]
  wire  m_175_io_x2; // @[MUL.scala 102:19]
  wire  m_175_io_x3; // @[MUL.scala 102:19]
  wire  m_175_io_s; // @[MUL.scala 102:19]
  wire  m_175_io_cout; // @[MUL.scala 102:19]
  wire  m_176_io_x1; // @[MUL.scala 102:19]
  wire  m_176_io_x2; // @[MUL.scala 102:19]
  wire  m_176_io_x3; // @[MUL.scala 102:19]
  wire  m_176_io_s; // @[MUL.scala 102:19]
  wire  m_176_io_cout; // @[MUL.scala 102:19]
  wire  m_177_io_x1; // @[MUL.scala 102:19]
  wire  m_177_io_x2; // @[MUL.scala 102:19]
  wire  m_177_io_x3; // @[MUL.scala 102:19]
  wire  m_177_io_s; // @[MUL.scala 102:19]
  wire  m_177_io_cout; // @[MUL.scala 102:19]
  wire  m_178_io_x1; // @[MUL.scala 102:19]
  wire  m_178_io_x2; // @[MUL.scala 102:19]
  wire  m_178_io_x3; // @[MUL.scala 102:19]
  wire  m_178_io_s; // @[MUL.scala 102:19]
  wire  m_178_io_cout; // @[MUL.scala 102:19]
  wire  m_179_io_x1; // @[MUL.scala 102:19]
  wire  m_179_io_x2; // @[MUL.scala 102:19]
  wire  m_179_io_x3; // @[MUL.scala 102:19]
  wire  m_179_io_s; // @[MUL.scala 102:19]
  wire  m_179_io_cout; // @[MUL.scala 102:19]
  wire  m_180_io_x1; // @[MUL.scala 102:19]
  wire  m_180_io_x2; // @[MUL.scala 102:19]
  wire  m_180_io_x3; // @[MUL.scala 102:19]
  wire  m_180_io_s; // @[MUL.scala 102:19]
  wire  m_180_io_cout; // @[MUL.scala 102:19]
  wire  m_181_io_x1; // @[MUL.scala 102:19]
  wire  m_181_io_x2; // @[MUL.scala 102:19]
  wire  m_181_io_x3; // @[MUL.scala 102:19]
  wire  m_181_io_s; // @[MUL.scala 102:19]
  wire  m_181_io_cout; // @[MUL.scala 102:19]
  wire  m_182_io_x1; // @[MUL.scala 102:19]
  wire  m_182_io_x2; // @[MUL.scala 102:19]
  wire  m_182_io_x3; // @[MUL.scala 102:19]
  wire  m_182_io_s; // @[MUL.scala 102:19]
  wire  m_182_io_cout; // @[MUL.scala 102:19]
  wire  m_183_io_x1; // @[MUL.scala 102:19]
  wire  m_183_io_x2; // @[MUL.scala 102:19]
  wire  m_183_io_x3; // @[MUL.scala 102:19]
  wire  m_183_io_s; // @[MUL.scala 102:19]
  wire  m_183_io_cout; // @[MUL.scala 102:19]
  wire  m_184_io_x1; // @[MUL.scala 102:19]
  wire  m_184_io_x2; // @[MUL.scala 102:19]
  wire  m_184_io_x3; // @[MUL.scala 102:19]
  wire  m_184_io_s; // @[MUL.scala 102:19]
  wire  m_184_io_cout; // @[MUL.scala 102:19]
  wire  m_185_io_x1; // @[MUL.scala 102:19]
  wire  m_185_io_x2; // @[MUL.scala 102:19]
  wire  m_185_io_x3; // @[MUL.scala 102:19]
  wire  m_185_io_s; // @[MUL.scala 102:19]
  wire  m_185_io_cout; // @[MUL.scala 102:19]
  wire  m_186_io_x1; // @[MUL.scala 102:19]
  wire  m_186_io_x2; // @[MUL.scala 102:19]
  wire  m_186_io_x3; // @[MUL.scala 102:19]
  wire  m_186_io_s; // @[MUL.scala 102:19]
  wire  m_186_io_cout; // @[MUL.scala 102:19]
  wire  m_187_io_x1; // @[MUL.scala 102:19]
  wire  m_187_io_x2; // @[MUL.scala 102:19]
  wire  m_187_io_x3; // @[MUL.scala 102:19]
  wire  m_187_io_s; // @[MUL.scala 102:19]
  wire  m_187_io_cout; // @[MUL.scala 102:19]
  wire  m_188_io_x1; // @[MUL.scala 102:19]
  wire  m_188_io_x2; // @[MUL.scala 102:19]
  wire  m_188_io_x3; // @[MUL.scala 102:19]
  wire  m_188_io_s; // @[MUL.scala 102:19]
  wire  m_188_io_cout; // @[MUL.scala 102:19]
  wire  m_189_io_x1; // @[MUL.scala 102:19]
  wire  m_189_io_x2; // @[MUL.scala 102:19]
  wire  m_189_io_x3; // @[MUL.scala 102:19]
  wire  m_189_io_s; // @[MUL.scala 102:19]
  wire  m_189_io_cout; // @[MUL.scala 102:19]
  wire  m_190_io_x1; // @[MUL.scala 102:19]
  wire  m_190_io_x2; // @[MUL.scala 102:19]
  wire  m_190_io_x3; // @[MUL.scala 102:19]
  wire  m_190_io_s; // @[MUL.scala 102:19]
  wire  m_190_io_cout; // @[MUL.scala 102:19]
  wire  m_191_io_x1; // @[MUL.scala 102:19]
  wire  m_191_io_x2; // @[MUL.scala 102:19]
  wire  m_191_io_x3; // @[MUL.scala 102:19]
  wire  m_191_io_s; // @[MUL.scala 102:19]
  wire  m_191_io_cout; // @[MUL.scala 102:19]
  wire  m_192_io_x1; // @[MUL.scala 102:19]
  wire  m_192_io_x2; // @[MUL.scala 102:19]
  wire  m_192_io_x3; // @[MUL.scala 102:19]
  wire  m_192_io_s; // @[MUL.scala 102:19]
  wire  m_192_io_cout; // @[MUL.scala 102:19]
  wire  m_193_io_in_0; // @[MUL.scala 124:19]
  wire  m_193_io_in_1; // @[MUL.scala 124:19]
  wire  m_193_io_out_0; // @[MUL.scala 124:19]
  wire  m_193_io_out_1; // @[MUL.scala 124:19]
  wire  m_194_io_x1; // @[MUL.scala 102:19]
  wire  m_194_io_x2; // @[MUL.scala 102:19]
  wire  m_194_io_x3; // @[MUL.scala 102:19]
  wire  m_194_io_s; // @[MUL.scala 102:19]
  wire  m_194_io_cout; // @[MUL.scala 102:19]
  wire  m_195_io_x1; // @[MUL.scala 102:19]
  wire  m_195_io_x2; // @[MUL.scala 102:19]
  wire  m_195_io_x3; // @[MUL.scala 102:19]
  wire  m_195_io_s; // @[MUL.scala 102:19]
  wire  m_195_io_cout; // @[MUL.scala 102:19]
  wire  m_196_io_x1; // @[MUL.scala 102:19]
  wire  m_196_io_x2; // @[MUL.scala 102:19]
  wire  m_196_io_x3; // @[MUL.scala 102:19]
  wire  m_196_io_s; // @[MUL.scala 102:19]
  wire  m_196_io_cout; // @[MUL.scala 102:19]
  wire  m_197_io_in_0; // @[MUL.scala 124:19]
  wire  m_197_io_in_1; // @[MUL.scala 124:19]
  wire  m_197_io_out_0; // @[MUL.scala 124:19]
  wire  m_197_io_out_1; // @[MUL.scala 124:19]
  wire  m_198_io_x1; // @[MUL.scala 102:19]
  wire  m_198_io_x2; // @[MUL.scala 102:19]
  wire  m_198_io_x3; // @[MUL.scala 102:19]
  wire  m_198_io_s; // @[MUL.scala 102:19]
  wire  m_198_io_cout; // @[MUL.scala 102:19]
  wire  m_199_io_x1; // @[MUL.scala 102:19]
  wire  m_199_io_x2; // @[MUL.scala 102:19]
  wire  m_199_io_x3; // @[MUL.scala 102:19]
  wire  m_199_io_s; // @[MUL.scala 102:19]
  wire  m_199_io_cout; // @[MUL.scala 102:19]
  wire  m_200_io_x1; // @[MUL.scala 102:19]
  wire  m_200_io_x2; // @[MUL.scala 102:19]
  wire  m_200_io_x3; // @[MUL.scala 102:19]
  wire  m_200_io_s; // @[MUL.scala 102:19]
  wire  m_200_io_cout; // @[MUL.scala 102:19]
  wire  m_201_io_x1; // @[MUL.scala 102:19]
  wire  m_201_io_x2; // @[MUL.scala 102:19]
  wire  m_201_io_x3; // @[MUL.scala 102:19]
  wire  m_201_io_s; // @[MUL.scala 102:19]
  wire  m_201_io_cout; // @[MUL.scala 102:19]
  wire  m_202_io_x1; // @[MUL.scala 102:19]
  wire  m_202_io_x2; // @[MUL.scala 102:19]
  wire  m_202_io_x3; // @[MUL.scala 102:19]
  wire  m_202_io_s; // @[MUL.scala 102:19]
  wire  m_202_io_cout; // @[MUL.scala 102:19]
  wire  m_203_io_x1; // @[MUL.scala 102:19]
  wire  m_203_io_x2; // @[MUL.scala 102:19]
  wire  m_203_io_x3; // @[MUL.scala 102:19]
  wire  m_203_io_s; // @[MUL.scala 102:19]
  wire  m_203_io_cout; // @[MUL.scala 102:19]
  wire  m_204_io_x1; // @[MUL.scala 102:19]
  wire  m_204_io_x2; // @[MUL.scala 102:19]
  wire  m_204_io_x3; // @[MUL.scala 102:19]
  wire  m_204_io_s; // @[MUL.scala 102:19]
  wire  m_204_io_cout; // @[MUL.scala 102:19]
  wire  m_205_io_x1; // @[MUL.scala 102:19]
  wire  m_205_io_x2; // @[MUL.scala 102:19]
  wire  m_205_io_x3; // @[MUL.scala 102:19]
  wire  m_205_io_s; // @[MUL.scala 102:19]
  wire  m_205_io_cout; // @[MUL.scala 102:19]
  wire  m_206_io_x1; // @[MUL.scala 102:19]
  wire  m_206_io_x2; // @[MUL.scala 102:19]
  wire  m_206_io_x3; // @[MUL.scala 102:19]
  wire  m_206_io_s; // @[MUL.scala 102:19]
  wire  m_206_io_cout; // @[MUL.scala 102:19]
  wire  m_207_io_x1; // @[MUL.scala 102:19]
  wire  m_207_io_x2; // @[MUL.scala 102:19]
  wire  m_207_io_x3; // @[MUL.scala 102:19]
  wire  m_207_io_s; // @[MUL.scala 102:19]
  wire  m_207_io_cout; // @[MUL.scala 102:19]
  wire  m_208_io_x1; // @[MUL.scala 102:19]
  wire  m_208_io_x2; // @[MUL.scala 102:19]
  wire  m_208_io_x3; // @[MUL.scala 102:19]
  wire  m_208_io_s; // @[MUL.scala 102:19]
  wire  m_208_io_cout; // @[MUL.scala 102:19]
  wire  m_209_io_x1; // @[MUL.scala 102:19]
  wire  m_209_io_x2; // @[MUL.scala 102:19]
  wire  m_209_io_x3; // @[MUL.scala 102:19]
  wire  m_209_io_s; // @[MUL.scala 102:19]
  wire  m_209_io_cout; // @[MUL.scala 102:19]
  wire  m_210_io_x1; // @[MUL.scala 102:19]
  wire  m_210_io_x2; // @[MUL.scala 102:19]
  wire  m_210_io_x3; // @[MUL.scala 102:19]
  wire  m_210_io_s; // @[MUL.scala 102:19]
  wire  m_210_io_cout; // @[MUL.scala 102:19]
  wire  m_211_io_x1; // @[MUL.scala 102:19]
  wire  m_211_io_x2; // @[MUL.scala 102:19]
  wire  m_211_io_x3; // @[MUL.scala 102:19]
  wire  m_211_io_s; // @[MUL.scala 102:19]
  wire  m_211_io_cout; // @[MUL.scala 102:19]
  wire  m_212_io_in_0; // @[MUL.scala 124:19]
  wire  m_212_io_in_1; // @[MUL.scala 124:19]
  wire  m_212_io_out_0; // @[MUL.scala 124:19]
  wire  m_212_io_out_1; // @[MUL.scala 124:19]
  wire  m_213_io_x1; // @[MUL.scala 102:19]
  wire  m_213_io_x2; // @[MUL.scala 102:19]
  wire  m_213_io_x3; // @[MUL.scala 102:19]
  wire  m_213_io_s; // @[MUL.scala 102:19]
  wire  m_213_io_cout; // @[MUL.scala 102:19]
  wire  m_214_io_x1; // @[MUL.scala 102:19]
  wire  m_214_io_x2; // @[MUL.scala 102:19]
  wire  m_214_io_x3; // @[MUL.scala 102:19]
  wire  m_214_io_s; // @[MUL.scala 102:19]
  wire  m_214_io_cout; // @[MUL.scala 102:19]
  wire  m_215_io_in_0; // @[MUL.scala 124:19]
  wire  m_215_io_in_1; // @[MUL.scala 124:19]
  wire  m_215_io_out_0; // @[MUL.scala 124:19]
  wire  m_215_io_out_1; // @[MUL.scala 124:19]
  wire  m_216_io_x1; // @[MUL.scala 102:19]
  wire  m_216_io_x2; // @[MUL.scala 102:19]
  wire  m_216_io_x3; // @[MUL.scala 102:19]
  wire  m_216_io_s; // @[MUL.scala 102:19]
  wire  m_216_io_cout; // @[MUL.scala 102:19]
  wire  m_217_io_x1; // @[MUL.scala 102:19]
  wire  m_217_io_x2; // @[MUL.scala 102:19]
  wire  m_217_io_x3; // @[MUL.scala 102:19]
  wire  m_217_io_s; // @[MUL.scala 102:19]
  wire  m_217_io_cout; // @[MUL.scala 102:19]
  wire  m_218_io_x1; // @[MUL.scala 102:19]
  wire  m_218_io_x2; // @[MUL.scala 102:19]
  wire  m_218_io_x3; // @[MUL.scala 102:19]
  wire  m_218_io_s; // @[MUL.scala 102:19]
  wire  m_218_io_cout; // @[MUL.scala 102:19]
  wire  m_219_io_x1; // @[MUL.scala 102:19]
  wire  m_219_io_x2; // @[MUL.scala 102:19]
  wire  m_219_io_x3; // @[MUL.scala 102:19]
  wire  m_219_io_s; // @[MUL.scala 102:19]
  wire  m_219_io_cout; // @[MUL.scala 102:19]
  wire  m_220_io_x1; // @[MUL.scala 102:19]
  wire  m_220_io_x2; // @[MUL.scala 102:19]
  wire  m_220_io_x3; // @[MUL.scala 102:19]
  wire  m_220_io_s; // @[MUL.scala 102:19]
  wire  m_220_io_cout; // @[MUL.scala 102:19]
  wire  m_221_io_x1; // @[MUL.scala 102:19]
  wire  m_221_io_x2; // @[MUL.scala 102:19]
  wire  m_221_io_x3; // @[MUL.scala 102:19]
  wire  m_221_io_s; // @[MUL.scala 102:19]
  wire  m_221_io_cout; // @[MUL.scala 102:19]
  wire  m_222_io_x1; // @[MUL.scala 102:19]
  wire  m_222_io_x2; // @[MUL.scala 102:19]
  wire  m_222_io_x3; // @[MUL.scala 102:19]
  wire  m_222_io_s; // @[MUL.scala 102:19]
  wire  m_222_io_cout; // @[MUL.scala 102:19]
  wire  m_223_io_x1; // @[MUL.scala 102:19]
  wire  m_223_io_x2; // @[MUL.scala 102:19]
  wire  m_223_io_x3; // @[MUL.scala 102:19]
  wire  m_223_io_s; // @[MUL.scala 102:19]
  wire  m_223_io_cout; // @[MUL.scala 102:19]
  wire  m_224_io_x1; // @[MUL.scala 102:19]
  wire  m_224_io_x2; // @[MUL.scala 102:19]
  wire  m_224_io_x3; // @[MUL.scala 102:19]
  wire  m_224_io_s; // @[MUL.scala 102:19]
  wire  m_224_io_cout; // @[MUL.scala 102:19]
  wire  m_225_io_in_0; // @[MUL.scala 124:19]
  wire  m_225_io_in_1; // @[MUL.scala 124:19]
  wire  m_225_io_out_0; // @[MUL.scala 124:19]
  wire  m_225_io_out_1; // @[MUL.scala 124:19]
  wire  m_226_io_x1; // @[MUL.scala 102:19]
  wire  m_226_io_x2; // @[MUL.scala 102:19]
  wire  m_226_io_x3; // @[MUL.scala 102:19]
  wire  m_226_io_s; // @[MUL.scala 102:19]
  wire  m_226_io_cout; // @[MUL.scala 102:19]
  wire  m_227_io_in_0; // @[MUL.scala 124:19]
  wire  m_227_io_in_1; // @[MUL.scala 124:19]
  wire  m_227_io_out_0; // @[MUL.scala 124:19]
  wire  m_227_io_out_1; // @[MUL.scala 124:19]
  wire  m_228_io_x1; // @[MUL.scala 102:19]
  wire  m_228_io_x2; // @[MUL.scala 102:19]
  wire  m_228_io_x3; // @[MUL.scala 102:19]
  wire  m_228_io_s; // @[MUL.scala 102:19]
  wire  m_228_io_cout; // @[MUL.scala 102:19]
  wire  m_229_io_x1; // @[MUL.scala 102:19]
  wire  m_229_io_x2; // @[MUL.scala 102:19]
  wire  m_229_io_x3; // @[MUL.scala 102:19]
  wire  m_229_io_s; // @[MUL.scala 102:19]
  wire  m_229_io_cout; // @[MUL.scala 102:19]
  wire  m_230_io_x1; // @[MUL.scala 102:19]
  wire  m_230_io_x2; // @[MUL.scala 102:19]
  wire  m_230_io_x3; // @[MUL.scala 102:19]
  wire  m_230_io_s; // @[MUL.scala 102:19]
  wire  m_230_io_cout; // @[MUL.scala 102:19]
  wire  m_231_io_x1; // @[MUL.scala 102:19]
  wire  m_231_io_x2; // @[MUL.scala 102:19]
  wire  m_231_io_x3; // @[MUL.scala 102:19]
  wire  m_231_io_s; // @[MUL.scala 102:19]
  wire  m_231_io_cout; // @[MUL.scala 102:19]
  wire  m_232_io_in_0; // @[MUL.scala 124:19]
  wire  m_232_io_in_1; // @[MUL.scala 124:19]
  wire  m_232_io_out_0; // @[MUL.scala 124:19]
  wire  m_232_io_out_1; // @[MUL.scala 124:19]
  wire  m_233_io_in_0; // @[MUL.scala 124:19]
  wire  m_233_io_in_1; // @[MUL.scala 124:19]
  wire  m_233_io_out_0; // @[MUL.scala 124:19]
  wire  m_233_io_out_1; // @[MUL.scala 124:19]
  wire  m_234_io_in_0; // @[MUL.scala 124:19]
  wire  m_234_io_in_1; // @[MUL.scala 124:19]
  wire  m_234_io_out_0; // @[MUL.scala 124:19]
  wire  m_234_io_out_1; // @[MUL.scala 124:19]
  wire  m_235_io_in_0; // @[MUL.scala 124:19]
  wire  m_235_io_in_1; // @[MUL.scala 124:19]
  wire  m_235_io_out_0; // @[MUL.scala 124:19]
  wire  m_235_io_out_1; // @[MUL.scala 124:19]
  wire  m_236_io_in_0; // @[MUL.scala 124:19]
  wire  m_236_io_in_1; // @[MUL.scala 124:19]
  wire  m_236_io_out_0; // @[MUL.scala 124:19]
  wire  m_236_io_out_1; // @[MUL.scala 124:19]
  wire  m_237_io_x1; // @[MUL.scala 102:19]
  wire  m_237_io_x2; // @[MUL.scala 102:19]
  wire  m_237_io_x3; // @[MUL.scala 102:19]
  wire  m_237_io_s; // @[MUL.scala 102:19]
  wire  m_237_io_cout; // @[MUL.scala 102:19]
  wire  m_238_io_x1; // @[MUL.scala 102:19]
  wire  m_238_io_x2; // @[MUL.scala 102:19]
  wire  m_238_io_x3; // @[MUL.scala 102:19]
  wire  m_238_io_s; // @[MUL.scala 102:19]
  wire  m_238_io_cout; // @[MUL.scala 102:19]
  wire  m_239_io_x1; // @[MUL.scala 102:19]
  wire  m_239_io_x2; // @[MUL.scala 102:19]
  wire  m_239_io_x3; // @[MUL.scala 102:19]
  wire  m_239_io_s; // @[MUL.scala 102:19]
  wire  m_239_io_cout; // @[MUL.scala 102:19]
  wire  m_240_io_x1; // @[MUL.scala 102:19]
  wire  m_240_io_x2; // @[MUL.scala 102:19]
  wire  m_240_io_x3; // @[MUL.scala 102:19]
  wire  m_240_io_s; // @[MUL.scala 102:19]
  wire  m_240_io_cout; // @[MUL.scala 102:19]
  wire  m_241_io_x1; // @[MUL.scala 102:19]
  wire  m_241_io_x2; // @[MUL.scala 102:19]
  wire  m_241_io_x3; // @[MUL.scala 102:19]
  wire  m_241_io_s; // @[MUL.scala 102:19]
  wire  m_241_io_cout; // @[MUL.scala 102:19]
  wire  m_242_io_x1; // @[MUL.scala 102:19]
  wire  m_242_io_x2; // @[MUL.scala 102:19]
  wire  m_242_io_x3; // @[MUL.scala 102:19]
  wire  m_242_io_s; // @[MUL.scala 102:19]
  wire  m_242_io_cout; // @[MUL.scala 102:19]
  wire  m_243_io_x1; // @[MUL.scala 102:19]
  wire  m_243_io_x2; // @[MUL.scala 102:19]
  wire  m_243_io_x3; // @[MUL.scala 102:19]
  wire  m_243_io_s; // @[MUL.scala 102:19]
  wire  m_243_io_cout; // @[MUL.scala 102:19]
  wire  m_244_io_in_0; // @[MUL.scala 124:19]
  wire  m_244_io_in_1; // @[MUL.scala 124:19]
  wire  m_244_io_out_0; // @[MUL.scala 124:19]
  wire  m_244_io_out_1; // @[MUL.scala 124:19]
  wire  m_245_io_x1; // @[MUL.scala 102:19]
  wire  m_245_io_x2; // @[MUL.scala 102:19]
  wire  m_245_io_x3; // @[MUL.scala 102:19]
  wire  m_245_io_s; // @[MUL.scala 102:19]
  wire  m_245_io_cout; // @[MUL.scala 102:19]
  wire  m_246_io_in_0; // @[MUL.scala 124:19]
  wire  m_246_io_in_1; // @[MUL.scala 124:19]
  wire  m_246_io_out_0; // @[MUL.scala 124:19]
  wire  m_246_io_out_1; // @[MUL.scala 124:19]
  wire  m_247_io_x1; // @[MUL.scala 102:19]
  wire  m_247_io_x2; // @[MUL.scala 102:19]
  wire  m_247_io_x3; // @[MUL.scala 102:19]
  wire  m_247_io_s; // @[MUL.scala 102:19]
  wire  m_247_io_cout; // @[MUL.scala 102:19]
  wire  m_248_io_in_0; // @[MUL.scala 124:19]
  wire  m_248_io_in_1; // @[MUL.scala 124:19]
  wire  m_248_io_out_0; // @[MUL.scala 124:19]
  wire  m_248_io_out_1; // @[MUL.scala 124:19]
  wire  m_249_io_x1; // @[MUL.scala 102:19]
  wire  m_249_io_x2; // @[MUL.scala 102:19]
  wire  m_249_io_x3; // @[MUL.scala 102:19]
  wire  m_249_io_s; // @[MUL.scala 102:19]
  wire  m_249_io_cout; // @[MUL.scala 102:19]
  wire  m_250_io_x1; // @[MUL.scala 102:19]
  wire  m_250_io_x2; // @[MUL.scala 102:19]
  wire  m_250_io_x3; // @[MUL.scala 102:19]
  wire  m_250_io_s; // @[MUL.scala 102:19]
  wire  m_250_io_cout; // @[MUL.scala 102:19]
  wire  m_251_io_x1; // @[MUL.scala 102:19]
  wire  m_251_io_x2; // @[MUL.scala 102:19]
  wire  m_251_io_x3; // @[MUL.scala 102:19]
  wire  m_251_io_s; // @[MUL.scala 102:19]
  wire  m_251_io_cout; // @[MUL.scala 102:19]
  wire  m_252_io_x1; // @[MUL.scala 102:19]
  wire  m_252_io_x2; // @[MUL.scala 102:19]
  wire  m_252_io_x3; // @[MUL.scala 102:19]
  wire  m_252_io_s; // @[MUL.scala 102:19]
  wire  m_252_io_cout; // @[MUL.scala 102:19]
  wire  m_253_io_x1; // @[MUL.scala 102:19]
  wire  m_253_io_x2; // @[MUL.scala 102:19]
  wire  m_253_io_x3; // @[MUL.scala 102:19]
  wire  m_253_io_s; // @[MUL.scala 102:19]
  wire  m_253_io_cout; // @[MUL.scala 102:19]
  wire  m_254_io_x1; // @[MUL.scala 102:19]
  wire  m_254_io_x2; // @[MUL.scala 102:19]
  wire  m_254_io_x3; // @[MUL.scala 102:19]
  wire  m_254_io_s; // @[MUL.scala 102:19]
  wire  m_254_io_cout; // @[MUL.scala 102:19]
  wire  m_255_io_x1; // @[MUL.scala 102:19]
  wire  m_255_io_x2; // @[MUL.scala 102:19]
  wire  m_255_io_x3; // @[MUL.scala 102:19]
  wire  m_255_io_s; // @[MUL.scala 102:19]
  wire  m_255_io_cout; // @[MUL.scala 102:19]
  wire  m_256_io_x1; // @[MUL.scala 102:19]
  wire  m_256_io_x2; // @[MUL.scala 102:19]
  wire  m_256_io_x3; // @[MUL.scala 102:19]
  wire  m_256_io_s; // @[MUL.scala 102:19]
  wire  m_256_io_cout; // @[MUL.scala 102:19]
  wire  m_257_io_x1; // @[MUL.scala 102:19]
  wire  m_257_io_x2; // @[MUL.scala 102:19]
  wire  m_257_io_x3; // @[MUL.scala 102:19]
  wire  m_257_io_s; // @[MUL.scala 102:19]
  wire  m_257_io_cout; // @[MUL.scala 102:19]
  wire  m_258_io_x1; // @[MUL.scala 102:19]
  wire  m_258_io_x2; // @[MUL.scala 102:19]
  wire  m_258_io_x3; // @[MUL.scala 102:19]
  wire  m_258_io_s; // @[MUL.scala 102:19]
  wire  m_258_io_cout; // @[MUL.scala 102:19]
  wire  m_259_io_x1; // @[MUL.scala 102:19]
  wire  m_259_io_x2; // @[MUL.scala 102:19]
  wire  m_259_io_x3; // @[MUL.scala 102:19]
  wire  m_259_io_s; // @[MUL.scala 102:19]
  wire  m_259_io_cout; // @[MUL.scala 102:19]
  wire  m_260_io_x1; // @[MUL.scala 102:19]
  wire  m_260_io_x2; // @[MUL.scala 102:19]
  wire  m_260_io_x3; // @[MUL.scala 102:19]
  wire  m_260_io_s; // @[MUL.scala 102:19]
  wire  m_260_io_cout; // @[MUL.scala 102:19]
  wire  m_261_io_x1; // @[MUL.scala 102:19]
  wire  m_261_io_x2; // @[MUL.scala 102:19]
  wire  m_261_io_x3; // @[MUL.scala 102:19]
  wire  m_261_io_s; // @[MUL.scala 102:19]
  wire  m_261_io_cout; // @[MUL.scala 102:19]
  wire  m_262_io_x1; // @[MUL.scala 102:19]
  wire  m_262_io_x2; // @[MUL.scala 102:19]
  wire  m_262_io_x3; // @[MUL.scala 102:19]
  wire  m_262_io_s; // @[MUL.scala 102:19]
  wire  m_262_io_cout; // @[MUL.scala 102:19]
  wire  m_263_io_in_0; // @[MUL.scala 124:19]
  wire  m_263_io_in_1; // @[MUL.scala 124:19]
  wire  m_263_io_out_0; // @[MUL.scala 124:19]
  wire  m_263_io_out_1; // @[MUL.scala 124:19]
  wire  m_264_io_x1; // @[MUL.scala 102:19]
  wire  m_264_io_x2; // @[MUL.scala 102:19]
  wire  m_264_io_x3; // @[MUL.scala 102:19]
  wire  m_264_io_s; // @[MUL.scala 102:19]
  wire  m_264_io_cout; // @[MUL.scala 102:19]
  wire  m_265_io_x1; // @[MUL.scala 102:19]
  wire  m_265_io_x2; // @[MUL.scala 102:19]
  wire  m_265_io_x3; // @[MUL.scala 102:19]
  wire  m_265_io_s; // @[MUL.scala 102:19]
  wire  m_265_io_cout; // @[MUL.scala 102:19]
  wire  m_266_io_in_0; // @[MUL.scala 124:19]
  wire  m_266_io_in_1; // @[MUL.scala 124:19]
  wire  m_266_io_out_0; // @[MUL.scala 124:19]
  wire  m_266_io_out_1; // @[MUL.scala 124:19]
  wire  m_267_io_x1; // @[MUL.scala 102:19]
  wire  m_267_io_x2; // @[MUL.scala 102:19]
  wire  m_267_io_x3; // @[MUL.scala 102:19]
  wire  m_267_io_s; // @[MUL.scala 102:19]
  wire  m_267_io_cout; // @[MUL.scala 102:19]
  wire  m_268_io_x1; // @[MUL.scala 102:19]
  wire  m_268_io_x2; // @[MUL.scala 102:19]
  wire  m_268_io_x3; // @[MUL.scala 102:19]
  wire  m_268_io_s; // @[MUL.scala 102:19]
  wire  m_268_io_cout; // @[MUL.scala 102:19]
  wire  m_269_io_in_0; // @[MUL.scala 124:19]
  wire  m_269_io_in_1; // @[MUL.scala 124:19]
  wire  m_269_io_out_0; // @[MUL.scala 124:19]
  wire  m_269_io_out_1; // @[MUL.scala 124:19]
  wire  m_270_io_x1; // @[MUL.scala 102:19]
  wire  m_270_io_x2; // @[MUL.scala 102:19]
  wire  m_270_io_x3; // @[MUL.scala 102:19]
  wire  m_270_io_s; // @[MUL.scala 102:19]
  wire  m_270_io_cout; // @[MUL.scala 102:19]
  wire  m_271_io_x1; // @[MUL.scala 102:19]
  wire  m_271_io_x2; // @[MUL.scala 102:19]
  wire  m_271_io_x3; // @[MUL.scala 102:19]
  wire  m_271_io_s; // @[MUL.scala 102:19]
  wire  m_271_io_cout; // @[MUL.scala 102:19]
  wire  m_272_io_x1; // @[MUL.scala 102:19]
  wire  m_272_io_x2; // @[MUL.scala 102:19]
  wire  m_272_io_x3; // @[MUL.scala 102:19]
  wire  m_272_io_s; // @[MUL.scala 102:19]
  wire  m_272_io_cout; // @[MUL.scala 102:19]
  wire  m_273_io_x1; // @[MUL.scala 102:19]
  wire  m_273_io_x2; // @[MUL.scala 102:19]
  wire  m_273_io_x3; // @[MUL.scala 102:19]
  wire  m_273_io_s; // @[MUL.scala 102:19]
  wire  m_273_io_cout; // @[MUL.scala 102:19]
  wire  m_274_io_x1; // @[MUL.scala 102:19]
  wire  m_274_io_x2; // @[MUL.scala 102:19]
  wire  m_274_io_x3; // @[MUL.scala 102:19]
  wire  m_274_io_s; // @[MUL.scala 102:19]
  wire  m_274_io_cout; // @[MUL.scala 102:19]
  wire  m_275_io_x1; // @[MUL.scala 102:19]
  wire  m_275_io_x2; // @[MUL.scala 102:19]
  wire  m_275_io_x3; // @[MUL.scala 102:19]
  wire  m_275_io_s; // @[MUL.scala 102:19]
  wire  m_275_io_cout; // @[MUL.scala 102:19]
  wire  m_276_io_x1; // @[MUL.scala 102:19]
  wire  m_276_io_x2; // @[MUL.scala 102:19]
  wire  m_276_io_x3; // @[MUL.scala 102:19]
  wire  m_276_io_s; // @[MUL.scala 102:19]
  wire  m_276_io_cout; // @[MUL.scala 102:19]
  wire  m_277_io_x1; // @[MUL.scala 102:19]
  wire  m_277_io_x2; // @[MUL.scala 102:19]
  wire  m_277_io_x3; // @[MUL.scala 102:19]
  wire  m_277_io_s; // @[MUL.scala 102:19]
  wire  m_277_io_cout; // @[MUL.scala 102:19]
  wire  m_278_io_x1; // @[MUL.scala 102:19]
  wire  m_278_io_x2; // @[MUL.scala 102:19]
  wire  m_278_io_x3; // @[MUL.scala 102:19]
  wire  m_278_io_s; // @[MUL.scala 102:19]
  wire  m_278_io_cout; // @[MUL.scala 102:19]
  wire  m_279_io_x1; // @[MUL.scala 102:19]
  wire  m_279_io_x2; // @[MUL.scala 102:19]
  wire  m_279_io_x3; // @[MUL.scala 102:19]
  wire  m_279_io_s; // @[MUL.scala 102:19]
  wire  m_279_io_cout; // @[MUL.scala 102:19]
  wire  m_280_io_x1; // @[MUL.scala 102:19]
  wire  m_280_io_x2; // @[MUL.scala 102:19]
  wire  m_280_io_x3; // @[MUL.scala 102:19]
  wire  m_280_io_s; // @[MUL.scala 102:19]
  wire  m_280_io_cout; // @[MUL.scala 102:19]
  wire  m_281_io_x1; // @[MUL.scala 102:19]
  wire  m_281_io_x2; // @[MUL.scala 102:19]
  wire  m_281_io_x3; // @[MUL.scala 102:19]
  wire  m_281_io_s; // @[MUL.scala 102:19]
  wire  m_281_io_cout; // @[MUL.scala 102:19]
  wire  m_282_io_x1; // @[MUL.scala 102:19]
  wire  m_282_io_x2; // @[MUL.scala 102:19]
  wire  m_282_io_x3; // @[MUL.scala 102:19]
  wire  m_282_io_s; // @[MUL.scala 102:19]
  wire  m_282_io_cout; // @[MUL.scala 102:19]
  wire  m_283_io_x1; // @[MUL.scala 102:19]
  wire  m_283_io_x2; // @[MUL.scala 102:19]
  wire  m_283_io_x3; // @[MUL.scala 102:19]
  wire  m_283_io_s; // @[MUL.scala 102:19]
  wire  m_283_io_cout; // @[MUL.scala 102:19]
  wire  m_284_io_x1; // @[MUL.scala 102:19]
  wire  m_284_io_x2; // @[MUL.scala 102:19]
  wire  m_284_io_x3; // @[MUL.scala 102:19]
  wire  m_284_io_s; // @[MUL.scala 102:19]
  wire  m_284_io_cout; // @[MUL.scala 102:19]
  wire  m_285_io_x1; // @[MUL.scala 102:19]
  wire  m_285_io_x2; // @[MUL.scala 102:19]
  wire  m_285_io_x3; // @[MUL.scala 102:19]
  wire  m_285_io_s; // @[MUL.scala 102:19]
  wire  m_285_io_cout; // @[MUL.scala 102:19]
  wire  m_286_io_x1; // @[MUL.scala 102:19]
  wire  m_286_io_x2; // @[MUL.scala 102:19]
  wire  m_286_io_x3; // @[MUL.scala 102:19]
  wire  m_286_io_s; // @[MUL.scala 102:19]
  wire  m_286_io_cout; // @[MUL.scala 102:19]
  wire  m_287_io_x1; // @[MUL.scala 102:19]
  wire  m_287_io_x2; // @[MUL.scala 102:19]
  wire  m_287_io_x3; // @[MUL.scala 102:19]
  wire  m_287_io_s; // @[MUL.scala 102:19]
  wire  m_287_io_cout; // @[MUL.scala 102:19]
  wire  m_288_io_x1; // @[MUL.scala 102:19]
  wire  m_288_io_x2; // @[MUL.scala 102:19]
  wire  m_288_io_x3; // @[MUL.scala 102:19]
  wire  m_288_io_s; // @[MUL.scala 102:19]
  wire  m_288_io_cout; // @[MUL.scala 102:19]
  wire  m_289_io_x1; // @[MUL.scala 102:19]
  wire  m_289_io_x2; // @[MUL.scala 102:19]
  wire  m_289_io_x3; // @[MUL.scala 102:19]
  wire  m_289_io_s; // @[MUL.scala 102:19]
  wire  m_289_io_cout; // @[MUL.scala 102:19]
  wire  m_290_io_x1; // @[MUL.scala 102:19]
  wire  m_290_io_x2; // @[MUL.scala 102:19]
  wire  m_290_io_x3; // @[MUL.scala 102:19]
  wire  m_290_io_s; // @[MUL.scala 102:19]
  wire  m_290_io_cout; // @[MUL.scala 102:19]
  wire  m_291_io_in_0; // @[MUL.scala 124:19]
  wire  m_291_io_in_1; // @[MUL.scala 124:19]
  wire  m_291_io_out_0; // @[MUL.scala 124:19]
  wire  m_291_io_out_1; // @[MUL.scala 124:19]
  wire  m_292_io_x1; // @[MUL.scala 102:19]
  wire  m_292_io_x2; // @[MUL.scala 102:19]
  wire  m_292_io_x3; // @[MUL.scala 102:19]
  wire  m_292_io_s; // @[MUL.scala 102:19]
  wire  m_292_io_cout; // @[MUL.scala 102:19]
  wire  m_293_io_x1; // @[MUL.scala 102:19]
  wire  m_293_io_x2; // @[MUL.scala 102:19]
  wire  m_293_io_x3; // @[MUL.scala 102:19]
  wire  m_293_io_s; // @[MUL.scala 102:19]
  wire  m_293_io_cout; // @[MUL.scala 102:19]
  wire  m_294_io_x1; // @[MUL.scala 102:19]
  wire  m_294_io_x2; // @[MUL.scala 102:19]
  wire  m_294_io_x3; // @[MUL.scala 102:19]
  wire  m_294_io_s; // @[MUL.scala 102:19]
  wire  m_294_io_cout; // @[MUL.scala 102:19]
  wire  m_295_io_in_0; // @[MUL.scala 124:19]
  wire  m_295_io_in_1; // @[MUL.scala 124:19]
  wire  m_295_io_out_0; // @[MUL.scala 124:19]
  wire  m_295_io_out_1; // @[MUL.scala 124:19]
  wire  m_296_io_x1; // @[MUL.scala 102:19]
  wire  m_296_io_x2; // @[MUL.scala 102:19]
  wire  m_296_io_x3; // @[MUL.scala 102:19]
  wire  m_296_io_s; // @[MUL.scala 102:19]
  wire  m_296_io_cout; // @[MUL.scala 102:19]
  wire  m_297_io_x1; // @[MUL.scala 102:19]
  wire  m_297_io_x2; // @[MUL.scala 102:19]
  wire  m_297_io_x3; // @[MUL.scala 102:19]
  wire  m_297_io_s; // @[MUL.scala 102:19]
  wire  m_297_io_cout; // @[MUL.scala 102:19]
  wire  m_298_io_x1; // @[MUL.scala 102:19]
  wire  m_298_io_x2; // @[MUL.scala 102:19]
  wire  m_298_io_x3; // @[MUL.scala 102:19]
  wire  m_298_io_s; // @[MUL.scala 102:19]
  wire  m_298_io_cout; // @[MUL.scala 102:19]
  wire  m_299_io_in_0; // @[MUL.scala 124:19]
  wire  m_299_io_in_1; // @[MUL.scala 124:19]
  wire  m_299_io_out_0; // @[MUL.scala 124:19]
  wire  m_299_io_out_1; // @[MUL.scala 124:19]
  wire  m_300_io_x1; // @[MUL.scala 102:19]
  wire  m_300_io_x2; // @[MUL.scala 102:19]
  wire  m_300_io_x3; // @[MUL.scala 102:19]
  wire  m_300_io_s; // @[MUL.scala 102:19]
  wire  m_300_io_cout; // @[MUL.scala 102:19]
  wire  m_301_io_x1; // @[MUL.scala 102:19]
  wire  m_301_io_x2; // @[MUL.scala 102:19]
  wire  m_301_io_x3; // @[MUL.scala 102:19]
  wire  m_301_io_s; // @[MUL.scala 102:19]
  wire  m_301_io_cout; // @[MUL.scala 102:19]
  wire  m_302_io_x1; // @[MUL.scala 102:19]
  wire  m_302_io_x2; // @[MUL.scala 102:19]
  wire  m_302_io_x3; // @[MUL.scala 102:19]
  wire  m_302_io_s; // @[MUL.scala 102:19]
  wire  m_302_io_cout; // @[MUL.scala 102:19]
  wire  m_303_io_x1; // @[MUL.scala 102:19]
  wire  m_303_io_x2; // @[MUL.scala 102:19]
  wire  m_303_io_x3; // @[MUL.scala 102:19]
  wire  m_303_io_s; // @[MUL.scala 102:19]
  wire  m_303_io_cout; // @[MUL.scala 102:19]
  wire  m_304_io_x1; // @[MUL.scala 102:19]
  wire  m_304_io_x2; // @[MUL.scala 102:19]
  wire  m_304_io_x3; // @[MUL.scala 102:19]
  wire  m_304_io_s; // @[MUL.scala 102:19]
  wire  m_304_io_cout; // @[MUL.scala 102:19]
  wire  m_305_io_x1; // @[MUL.scala 102:19]
  wire  m_305_io_x2; // @[MUL.scala 102:19]
  wire  m_305_io_x3; // @[MUL.scala 102:19]
  wire  m_305_io_s; // @[MUL.scala 102:19]
  wire  m_305_io_cout; // @[MUL.scala 102:19]
  wire  m_306_io_x1; // @[MUL.scala 102:19]
  wire  m_306_io_x2; // @[MUL.scala 102:19]
  wire  m_306_io_x3; // @[MUL.scala 102:19]
  wire  m_306_io_s; // @[MUL.scala 102:19]
  wire  m_306_io_cout; // @[MUL.scala 102:19]
  wire  m_307_io_x1; // @[MUL.scala 102:19]
  wire  m_307_io_x2; // @[MUL.scala 102:19]
  wire  m_307_io_x3; // @[MUL.scala 102:19]
  wire  m_307_io_s; // @[MUL.scala 102:19]
  wire  m_307_io_cout; // @[MUL.scala 102:19]
  wire  m_308_io_x1; // @[MUL.scala 102:19]
  wire  m_308_io_x2; // @[MUL.scala 102:19]
  wire  m_308_io_x3; // @[MUL.scala 102:19]
  wire  m_308_io_s; // @[MUL.scala 102:19]
  wire  m_308_io_cout; // @[MUL.scala 102:19]
  wire  m_309_io_x1; // @[MUL.scala 102:19]
  wire  m_309_io_x2; // @[MUL.scala 102:19]
  wire  m_309_io_x3; // @[MUL.scala 102:19]
  wire  m_309_io_s; // @[MUL.scala 102:19]
  wire  m_309_io_cout; // @[MUL.scala 102:19]
  wire  m_310_io_x1; // @[MUL.scala 102:19]
  wire  m_310_io_x2; // @[MUL.scala 102:19]
  wire  m_310_io_x3; // @[MUL.scala 102:19]
  wire  m_310_io_s; // @[MUL.scala 102:19]
  wire  m_310_io_cout; // @[MUL.scala 102:19]
  wire  m_311_io_x1; // @[MUL.scala 102:19]
  wire  m_311_io_x2; // @[MUL.scala 102:19]
  wire  m_311_io_x3; // @[MUL.scala 102:19]
  wire  m_311_io_s; // @[MUL.scala 102:19]
  wire  m_311_io_cout; // @[MUL.scala 102:19]
  wire  m_312_io_x1; // @[MUL.scala 102:19]
  wire  m_312_io_x2; // @[MUL.scala 102:19]
  wire  m_312_io_x3; // @[MUL.scala 102:19]
  wire  m_312_io_s; // @[MUL.scala 102:19]
  wire  m_312_io_cout; // @[MUL.scala 102:19]
  wire  m_313_io_x1; // @[MUL.scala 102:19]
  wire  m_313_io_x2; // @[MUL.scala 102:19]
  wire  m_313_io_x3; // @[MUL.scala 102:19]
  wire  m_313_io_s; // @[MUL.scala 102:19]
  wire  m_313_io_cout; // @[MUL.scala 102:19]
  wire  m_314_io_x1; // @[MUL.scala 102:19]
  wire  m_314_io_x2; // @[MUL.scala 102:19]
  wire  m_314_io_x3; // @[MUL.scala 102:19]
  wire  m_314_io_s; // @[MUL.scala 102:19]
  wire  m_314_io_cout; // @[MUL.scala 102:19]
  wire  m_315_io_x1; // @[MUL.scala 102:19]
  wire  m_315_io_x2; // @[MUL.scala 102:19]
  wire  m_315_io_x3; // @[MUL.scala 102:19]
  wire  m_315_io_s; // @[MUL.scala 102:19]
  wire  m_315_io_cout; // @[MUL.scala 102:19]
  wire  m_316_io_x1; // @[MUL.scala 102:19]
  wire  m_316_io_x2; // @[MUL.scala 102:19]
  wire  m_316_io_x3; // @[MUL.scala 102:19]
  wire  m_316_io_s; // @[MUL.scala 102:19]
  wire  m_316_io_cout; // @[MUL.scala 102:19]
  wire  m_317_io_x1; // @[MUL.scala 102:19]
  wire  m_317_io_x2; // @[MUL.scala 102:19]
  wire  m_317_io_x3; // @[MUL.scala 102:19]
  wire  m_317_io_s; // @[MUL.scala 102:19]
  wire  m_317_io_cout; // @[MUL.scala 102:19]
  wire  m_318_io_x1; // @[MUL.scala 102:19]
  wire  m_318_io_x2; // @[MUL.scala 102:19]
  wire  m_318_io_x3; // @[MUL.scala 102:19]
  wire  m_318_io_s; // @[MUL.scala 102:19]
  wire  m_318_io_cout; // @[MUL.scala 102:19]
  wire  m_319_io_x1; // @[MUL.scala 102:19]
  wire  m_319_io_x2; // @[MUL.scala 102:19]
  wire  m_319_io_x3; // @[MUL.scala 102:19]
  wire  m_319_io_s; // @[MUL.scala 102:19]
  wire  m_319_io_cout; // @[MUL.scala 102:19]
  wire  m_320_io_x1; // @[MUL.scala 102:19]
  wire  m_320_io_x2; // @[MUL.scala 102:19]
  wire  m_320_io_x3; // @[MUL.scala 102:19]
  wire  m_320_io_s; // @[MUL.scala 102:19]
  wire  m_320_io_cout; // @[MUL.scala 102:19]
  wire  m_321_io_x1; // @[MUL.scala 102:19]
  wire  m_321_io_x2; // @[MUL.scala 102:19]
  wire  m_321_io_x3; // @[MUL.scala 102:19]
  wire  m_321_io_s; // @[MUL.scala 102:19]
  wire  m_321_io_cout; // @[MUL.scala 102:19]
  wire  m_322_io_x1; // @[MUL.scala 102:19]
  wire  m_322_io_x2; // @[MUL.scala 102:19]
  wire  m_322_io_x3; // @[MUL.scala 102:19]
  wire  m_322_io_s; // @[MUL.scala 102:19]
  wire  m_322_io_cout; // @[MUL.scala 102:19]
  wire  m_323_io_x1; // @[MUL.scala 102:19]
  wire  m_323_io_x2; // @[MUL.scala 102:19]
  wire  m_323_io_x3; // @[MUL.scala 102:19]
  wire  m_323_io_s; // @[MUL.scala 102:19]
  wire  m_323_io_cout; // @[MUL.scala 102:19]
  wire  m_324_io_x1; // @[MUL.scala 102:19]
  wire  m_324_io_x2; // @[MUL.scala 102:19]
  wire  m_324_io_x3; // @[MUL.scala 102:19]
  wire  m_324_io_s; // @[MUL.scala 102:19]
  wire  m_324_io_cout; // @[MUL.scala 102:19]
  wire  m_325_io_x1; // @[MUL.scala 102:19]
  wire  m_325_io_x2; // @[MUL.scala 102:19]
  wire  m_325_io_x3; // @[MUL.scala 102:19]
  wire  m_325_io_s; // @[MUL.scala 102:19]
  wire  m_325_io_cout; // @[MUL.scala 102:19]
  wire  m_326_io_x1; // @[MUL.scala 102:19]
  wire  m_326_io_x2; // @[MUL.scala 102:19]
  wire  m_326_io_x3; // @[MUL.scala 102:19]
  wire  m_326_io_s; // @[MUL.scala 102:19]
  wire  m_326_io_cout; // @[MUL.scala 102:19]
  wire  m_327_io_x1; // @[MUL.scala 102:19]
  wire  m_327_io_x2; // @[MUL.scala 102:19]
  wire  m_327_io_x3; // @[MUL.scala 102:19]
  wire  m_327_io_s; // @[MUL.scala 102:19]
  wire  m_327_io_cout; // @[MUL.scala 102:19]
  wire  m_328_io_x1; // @[MUL.scala 102:19]
  wire  m_328_io_x2; // @[MUL.scala 102:19]
  wire  m_328_io_x3; // @[MUL.scala 102:19]
  wire  m_328_io_s; // @[MUL.scala 102:19]
  wire  m_328_io_cout; // @[MUL.scala 102:19]
  wire  m_329_io_x1; // @[MUL.scala 102:19]
  wire  m_329_io_x2; // @[MUL.scala 102:19]
  wire  m_329_io_x3; // @[MUL.scala 102:19]
  wire  m_329_io_s; // @[MUL.scala 102:19]
  wire  m_329_io_cout; // @[MUL.scala 102:19]
  wire  m_330_io_x1; // @[MUL.scala 102:19]
  wire  m_330_io_x2; // @[MUL.scala 102:19]
  wire  m_330_io_x3; // @[MUL.scala 102:19]
  wire  m_330_io_s; // @[MUL.scala 102:19]
  wire  m_330_io_cout; // @[MUL.scala 102:19]
  wire  m_331_io_x1; // @[MUL.scala 102:19]
  wire  m_331_io_x2; // @[MUL.scala 102:19]
  wire  m_331_io_x3; // @[MUL.scala 102:19]
  wire  m_331_io_s; // @[MUL.scala 102:19]
  wire  m_331_io_cout; // @[MUL.scala 102:19]
  wire  m_332_io_x1; // @[MUL.scala 102:19]
  wire  m_332_io_x2; // @[MUL.scala 102:19]
  wire  m_332_io_x3; // @[MUL.scala 102:19]
  wire  m_332_io_s; // @[MUL.scala 102:19]
  wire  m_332_io_cout; // @[MUL.scala 102:19]
  wire  m_333_io_x1; // @[MUL.scala 102:19]
  wire  m_333_io_x2; // @[MUL.scala 102:19]
  wire  m_333_io_x3; // @[MUL.scala 102:19]
  wire  m_333_io_s; // @[MUL.scala 102:19]
  wire  m_333_io_cout; // @[MUL.scala 102:19]
  wire  m_334_io_x1; // @[MUL.scala 102:19]
  wire  m_334_io_x2; // @[MUL.scala 102:19]
  wire  m_334_io_x3; // @[MUL.scala 102:19]
  wire  m_334_io_s; // @[MUL.scala 102:19]
  wire  m_334_io_cout; // @[MUL.scala 102:19]
  wire  m_335_io_x1; // @[MUL.scala 102:19]
  wire  m_335_io_x2; // @[MUL.scala 102:19]
  wire  m_335_io_x3; // @[MUL.scala 102:19]
  wire  m_335_io_s; // @[MUL.scala 102:19]
  wire  m_335_io_cout; // @[MUL.scala 102:19]
  wire  m_336_io_x1; // @[MUL.scala 102:19]
  wire  m_336_io_x2; // @[MUL.scala 102:19]
  wire  m_336_io_x3; // @[MUL.scala 102:19]
  wire  m_336_io_s; // @[MUL.scala 102:19]
  wire  m_336_io_cout; // @[MUL.scala 102:19]
  wire  m_337_io_x1; // @[MUL.scala 102:19]
  wire  m_337_io_x2; // @[MUL.scala 102:19]
  wire  m_337_io_x3; // @[MUL.scala 102:19]
  wire  m_337_io_s; // @[MUL.scala 102:19]
  wire  m_337_io_cout; // @[MUL.scala 102:19]
  wire  m_338_io_x1; // @[MUL.scala 102:19]
  wire  m_338_io_x2; // @[MUL.scala 102:19]
  wire  m_338_io_x3; // @[MUL.scala 102:19]
  wire  m_338_io_s; // @[MUL.scala 102:19]
  wire  m_338_io_cout; // @[MUL.scala 102:19]
  wire  m_339_io_x1; // @[MUL.scala 102:19]
  wire  m_339_io_x2; // @[MUL.scala 102:19]
  wire  m_339_io_x3; // @[MUL.scala 102:19]
  wire  m_339_io_s; // @[MUL.scala 102:19]
  wire  m_339_io_cout; // @[MUL.scala 102:19]
  wire  m_340_io_x1; // @[MUL.scala 102:19]
  wire  m_340_io_x2; // @[MUL.scala 102:19]
  wire  m_340_io_x3; // @[MUL.scala 102:19]
  wire  m_340_io_s; // @[MUL.scala 102:19]
  wire  m_340_io_cout; // @[MUL.scala 102:19]
  wire  m_341_io_x1; // @[MUL.scala 102:19]
  wire  m_341_io_x2; // @[MUL.scala 102:19]
  wire  m_341_io_x3; // @[MUL.scala 102:19]
  wire  m_341_io_s; // @[MUL.scala 102:19]
  wire  m_341_io_cout; // @[MUL.scala 102:19]
  wire  m_342_io_x1; // @[MUL.scala 102:19]
  wire  m_342_io_x2; // @[MUL.scala 102:19]
  wire  m_342_io_x3; // @[MUL.scala 102:19]
  wire  m_342_io_s; // @[MUL.scala 102:19]
  wire  m_342_io_cout; // @[MUL.scala 102:19]
  wire  m_343_io_x1; // @[MUL.scala 102:19]
  wire  m_343_io_x2; // @[MUL.scala 102:19]
  wire  m_343_io_x3; // @[MUL.scala 102:19]
  wire  m_343_io_s; // @[MUL.scala 102:19]
  wire  m_343_io_cout; // @[MUL.scala 102:19]
  wire  m_344_io_x1; // @[MUL.scala 102:19]
  wire  m_344_io_x2; // @[MUL.scala 102:19]
  wire  m_344_io_x3; // @[MUL.scala 102:19]
  wire  m_344_io_s; // @[MUL.scala 102:19]
  wire  m_344_io_cout; // @[MUL.scala 102:19]
  wire  m_345_io_x1; // @[MUL.scala 102:19]
  wire  m_345_io_x2; // @[MUL.scala 102:19]
  wire  m_345_io_x3; // @[MUL.scala 102:19]
  wire  m_345_io_s; // @[MUL.scala 102:19]
  wire  m_345_io_cout; // @[MUL.scala 102:19]
  wire  m_346_io_x1; // @[MUL.scala 102:19]
  wire  m_346_io_x2; // @[MUL.scala 102:19]
  wire  m_346_io_x3; // @[MUL.scala 102:19]
  wire  m_346_io_s; // @[MUL.scala 102:19]
  wire  m_346_io_cout; // @[MUL.scala 102:19]
  wire  m_347_io_x1; // @[MUL.scala 102:19]
  wire  m_347_io_x2; // @[MUL.scala 102:19]
  wire  m_347_io_x3; // @[MUL.scala 102:19]
  wire  m_347_io_s; // @[MUL.scala 102:19]
  wire  m_347_io_cout; // @[MUL.scala 102:19]
  wire  m_348_io_in_0; // @[MUL.scala 124:19]
  wire  m_348_io_in_1; // @[MUL.scala 124:19]
  wire  m_348_io_out_0; // @[MUL.scala 124:19]
  wire  m_348_io_out_1; // @[MUL.scala 124:19]
  wire  m_349_io_x1; // @[MUL.scala 102:19]
  wire  m_349_io_x2; // @[MUL.scala 102:19]
  wire  m_349_io_x3; // @[MUL.scala 102:19]
  wire  m_349_io_s; // @[MUL.scala 102:19]
  wire  m_349_io_cout; // @[MUL.scala 102:19]
  wire  m_350_io_x1; // @[MUL.scala 102:19]
  wire  m_350_io_x2; // @[MUL.scala 102:19]
  wire  m_350_io_x3; // @[MUL.scala 102:19]
  wire  m_350_io_s; // @[MUL.scala 102:19]
  wire  m_350_io_cout; // @[MUL.scala 102:19]
  wire  m_351_io_in_0; // @[MUL.scala 124:19]
  wire  m_351_io_in_1; // @[MUL.scala 124:19]
  wire  m_351_io_out_0; // @[MUL.scala 124:19]
  wire  m_351_io_out_1; // @[MUL.scala 124:19]
  wire  m_352_io_x1; // @[MUL.scala 102:19]
  wire  m_352_io_x2; // @[MUL.scala 102:19]
  wire  m_352_io_x3; // @[MUL.scala 102:19]
  wire  m_352_io_s; // @[MUL.scala 102:19]
  wire  m_352_io_cout; // @[MUL.scala 102:19]
  wire  m_353_io_x1; // @[MUL.scala 102:19]
  wire  m_353_io_x2; // @[MUL.scala 102:19]
  wire  m_353_io_x3; // @[MUL.scala 102:19]
  wire  m_353_io_s; // @[MUL.scala 102:19]
  wire  m_353_io_cout; // @[MUL.scala 102:19]
  wire  m_354_io_in_0; // @[MUL.scala 124:19]
  wire  m_354_io_in_1; // @[MUL.scala 124:19]
  wire  m_354_io_out_0; // @[MUL.scala 124:19]
  wire  m_354_io_out_1; // @[MUL.scala 124:19]
  wire  m_355_io_x1; // @[MUL.scala 102:19]
  wire  m_355_io_x2; // @[MUL.scala 102:19]
  wire  m_355_io_x3; // @[MUL.scala 102:19]
  wire  m_355_io_s; // @[MUL.scala 102:19]
  wire  m_355_io_cout; // @[MUL.scala 102:19]
  wire  m_356_io_x1; // @[MUL.scala 102:19]
  wire  m_356_io_x2; // @[MUL.scala 102:19]
  wire  m_356_io_x3; // @[MUL.scala 102:19]
  wire  m_356_io_s; // @[MUL.scala 102:19]
  wire  m_356_io_cout; // @[MUL.scala 102:19]
  wire  m_357_io_in_0; // @[MUL.scala 124:19]
  wire  m_357_io_in_1; // @[MUL.scala 124:19]
  wire  m_357_io_out_0; // @[MUL.scala 124:19]
  wire  m_357_io_out_1; // @[MUL.scala 124:19]
  wire  m_358_io_x1; // @[MUL.scala 102:19]
  wire  m_358_io_x2; // @[MUL.scala 102:19]
  wire  m_358_io_x3; // @[MUL.scala 102:19]
  wire  m_358_io_s; // @[MUL.scala 102:19]
  wire  m_358_io_cout; // @[MUL.scala 102:19]
  wire  m_359_io_x1; // @[MUL.scala 102:19]
  wire  m_359_io_x2; // @[MUL.scala 102:19]
  wire  m_359_io_x3; // @[MUL.scala 102:19]
  wire  m_359_io_s; // @[MUL.scala 102:19]
  wire  m_359_io_cout; // @[MUL.scala 102:19]
  wire  m_360_io_in_0; // @[MUL.scala 124:19]
  wire  m_360_io_in_1; // @[MUL.scala 124:19]
  wire  m_360_io_out_0; // @[MUL.scala 124:19]
  wire  m_360_io_out_1; // @[MUL.scala 124:19]
  wire  m_361_io_x1; // @[MUL.scala 102:19]
  wire  m_361_io_x2; // @[MUL.scala 102:19]
  wire  m_361_io_x3; // @[MUL.scala 102:19]
  wire  m_361_io_s; // @[MUL.scala 102:19]
  wire  m_361_io_cout; // @[MUL.scala 102:19]
  wire  m_362_io_x1; // @[MUL.scala 102:19]
  wire  m_362_io_x2; // @[MUL.scala 102:19]
  wire  m_362_io_x3; // @[MUL.scala 102:19]
  wire  m_362_io_s; // @[MUL.scala 102:19]
  wire  m_362_io_cout; // @[MUL.scala 102:19]
  wire  m_363_io_x1; // @[MUL.scala 102:19]
  wire  m_363_io_x2; // @[MUL.scala 102:19]
  wire  m_363_io_x3; // @[MUL.scala 102:19]
  wire  m_363_io_s; // @[MUL.scala 102:19]
  wire  m_363_io_cout; // @[MUL.scala 102:19]
  wire  m_364_io_x1; // @[MUL.scala 102:19]
  wire  m_364_io_x2; // @[MUL.scala 102:19]
  wire  m_364_io_x3; // @[MUL.scala 102:19]
  wire  m_364_io_s; // @[MUL.scala 102:19]
  wire  m_364_io_cout; // @[MUL.scala 102:19]
  wire  m_365_io_x1; // @[MUL.scala 102:19]
  wire  m_365_io_x2; // @[MUL.scala 102:19]
  wire  m_365_io_x3; // @[MUL.scala 102:19]
  wire  m_365_io_s; // @[MUL.scala 102:19]
  wire  m_365_io_cout; // @[MUL.scala 102:19]
  wire  m_366_io_x1; // @[MUL.scala 102:19]
  wire  m_366_io_x2; // @[MUL.scala 102:19]
  wire  m_366_io_x3; // @[MUL.scala 102:19]
  wire  m_366_io_s; // @[MUL.scala 102:19]
  wire  m_366_io_cout; // @[MUL.scala 102:19]
  wire  m_367_io_x1; // @[MUL.scala 102:19]
  wire  m_367_io_x2; // @[MUL.scala 102:19]
  wire  m_367_io_x3; // @[MUL.scala 102:19]
  wire  m_367_io_s; // @[MUL.scala 102:19]
  wire  m_367_io_cout; // @[MUL.scala 102:19]
  wire  m_368_io_x1; // @[MUL.scala 102:19]
  wire  m_368_io_x2; // @[MUL.scala 102:19]
  wire  m_368_io_x3; // @[MUL.scala 102:19]
  wire  m_368_io_s; // @[MUL.scala 102:19]
  wire  m_368_io_cout; // @[MUL.scala 102:19]
  wire  m_369_io_x1; // @[MUL.scala 102:19]
  wire  m_369_io_x2; // @[MUL.scala 102:19]
  wire  m_369_io_x3; // @[MUL.scala 102:19]
  wire  m_369_io_s; // @[MUL.scala 102:19]
  wire  m_369_io_cout; // @[MUL.scala 102:19]
  wire  m_370_io_x1; // @[MUL.scala 102:19]
  wire  m_370_io_x2; // @[MUL.scala 102:19]
  wire  m_370_io_x3; // @[MUL.scala 102:19]
  wire  m_370_io_s; // @[MUL.scala 102:19]
  wire  m_370_io_cout; // @[MUL.scala 102:19]
  wire  m_371_io_x1; // @[MUL.scala 102:19]
  wire  m_371_io_x2; // @[MUL.scala 102:19]
  wire  m_371_io_x3; // @[MUL.scala 102:19]
  wire  m_371_io_s; // @[MUL.scala 102:19]
  wire  m_371_io_cout; // @[MUL.scala 102:19]
  wire  m_372_io_x1; // @[MUL.scala 102:19]
  wire  m_372_io_x2; // @[MUL.scala 102:19]
  wire  m_372_io_x3; // @[MUL.scala 102:19]
  wire  m_372_io_s; // @[MUL.scala 102:19]
  wire  m_372_io_cout; // @[MUL.scala 102:19]
  wire  m_373_io_x1; // @[MUL.scala 102:19]
  wire  m_373_io_x2; // @[MUL.scala 102:19]
  wire  m_373_io_x3; // @[MUL.scala 102:19]
  wire  m_373_io_s; // @[MUL.scala 102:19]
  wire  m_373_io_cout; // @[MUL.scala 102:19]
  wire  m_374_io_in_0; // @[MUL.scala 124:19]
  wire  m_374_io_in_1; // @[MUL.scala 124:19]
  wire  m_374_io_out_0; // @[MUL.scala 124:19]
  wire  m_374_io_out_1; // @[MUL.scala 124:19]
  wire  m_375_io_x1; // @[MUL.scala 102:19]
  wire  m_375_io_x2; // @[MUL.scala 102:19]
  wire  m_375_io_x3; // @[MUL.scala 102:19]
  wire  m_375_io_s; // @[MUL.scala 102:19]
  wire  m_375_io_cout; // @[MUL.scala 102:19]
  wire  m_376_io_x1; // @[MUL.scala 102:19]
  wire  m_376_io_x2; // @[MUL.scala 102:19]
  wire  m_376_io_x3; // @[MUL.scala 102:19]
  wire  m_376_io_s; // @[MUL.scala 102:19]
  wire  m_376_io_cout; // @[MUL.scala 102:19]
  wire  m_377_io_x1; // @[MUL.scala 102:19]
  wire  m_377_io_x2; // @[MUL.scala 102:19]
  wire  m_377_io_x3; // @[MUL.scala 102:19]
  wire  m_377_io_s; // @[MUL.scala 102:19]
  wire  m_377_io_cout; // @[MUL.scala 102:19]
  wire  m_378_io_x1; // @[MUL.scala 102:19]
  wire  m_378_io_x2; // @[MUL.scala 102:19]
  wire  m_378_io_x3; // @[MUL.scala 102:19]
  wire  m_378_io_s; // @[MUL.scala 102:19]
  wire  m_378_io_cout; // @[MUL.scala 102:19]
  wire  m_379_io_x1; // @[MUL.scala 102:19]
  wire  m_379_io_x2; // @[MUL.scala 102:19]
  wire  m_379_io_x3; // @[MUL.scala 102:19]
  wire  m_379_io_s; // @[MUL.scala 102:19]
  wire  m_379_io_cout; // @[MUL.scala 102:19]
  wire  m_380_io_x1; // @[MUL.scala 102:19]
  wire  m_380_io_x2; // @[MUL.scala 102:19]
  wire  m_380_io_x3; // @[MUL.scala 102:19]
  wire  m_380_io_s; // @[MUL.scala 102:19]
  wire  m_380_io_cout; // @[MUL.scala 102:19]
  wire  m_381_io_in_0; // @[MUL.scala 124:19]
  wire  m_381_io_in_1; // @[MUL.scala 124:19]
  wire  m_381_io_out_0; // @[MUL.scala 124:19]
  wire  m_381_io_out_1; // @[MUL.scala 124:19]
  wire  m_382_io_in_0; // @[MUL.scala 124:19]
  wire  m_382_io_in_1; // @[MUL.scala 124:19]
  wire  m_382_io_out_0; // @[MUL.scala 124:19]
  wire  m_382_io_out_1; // @[MUL.scala 124:19]
  wire  m_383_io_in_0; // @[MUL.scala 124:19]
  wire  m_383_io_in_1; // @[MUL.scala 124:19]
  wire  m_383_io_out_0; // @[MUL.scala 124:19]
  wire  m_383_io_out_1; // @[MUL.scala 124:19]
  wire  m_384_io_in_0; // @[MUL.scala 124:19]
  wire  m_384_io_in_1; // @[MUL.scala 124:19]
  wire  m_384_io_out_0; // @[MUL.scala 124:19]
  wire  m_384_io_out_1; // @[MUL.scala 124:19]
  wire  m_385_io_in_0; // @[MUL.scala 124:19]
  wire  m_385_io_in_1; // @[MUL.scala 124:19]
  wire  m_385_io_out_0; // @[MUL.scala 124:19]
  wire  m_385_io_out_1; // @[MUL.scala 124:19]
  wire  m_386_io_in_0; // @[MUL.scala 124:19]
  wire  m_386_io_in_1; // @[MUL.scala 124:19]
  wire  m_386_io_out_0; // @[MUL.scala 124:19]
  wire  m_386_io_out_1; // @[MUL.scala 124:19]
  wire  m_387_io_in_0; // @[MUL.scala 124:19]
  wire  m_387_io_in_1; // @[MUL.scala 124:19]
  wire  m_387_io_out_0; // @[MUL.scala 124:19]
  wire  m_387_io_out_1; // @[MUL.scala 124:19]
  wire  m_388_io_in_0; // @[MUL.scala 124:19]
  wire  m_388_io_in_1; // @[MUL.scala 124:19]
  wire  m_388_io_out_0; // @[MUL.scala 124:19]
  wire  m_388_io_out_1; // @[MUL.scala 124:19]
  wire  m_389_io_in_0; // @[MUL.scala 124:19]
  wire  m_389_io_in_1; // @[MUL.scala 124:19]
  wire  m_389_io_out_0; // @[MUL.scala 124:19]
  wire  m_389_io_out_1; // @[MUL.scala 124:19]
  wire  m_390_io_in_0; // @[MUL.scala 124:19]
  wire  m_390_io_in_1; // @[MUL.scala 124:19]
  wire  m_390_io_out_0; // @[MUL.scala 124:19]
  wire  m_390_io_out_1; // @[MUL.scala 124:19]
  wire  m_391_io_x1; // @[MUL.scala 102:19]
  wire  m_391_io_x2; // @[MUL.scala 102:19]
  wire  m_391_io_x3; // @[MUL.scala 102:19]
  wire  m_391_io_s; // @[MUL.scala 102:19]
  wire  m_391_io_cout; // @[MUL.scala 102:19]
  wire  m_392_io_x1; // @[MUL.scala 102:19]
  wire  m_392_io_x2; // @[MUL.scala 102:19]
  wire  m_392_io_x3; // @[MUL.scala 102:19]
  wire  m_392_io_s; // @[MUL.scala 102:19]
  wire  m_392_io_cout; // @[MUL.scala 102:19]
  wire  m_393_io_x1; // @[MUL.scala 102:19]
  wire  m_393_io_x2; // @[MUL.scala 102:19]
  wire  m_393_io_x3; // @[MUL.scala 102:19]
  wire  m_393_io_s; // @[MUL.scala 102:19]
  wire  m_393_io_cout; // @[MUL.scala 102:19]
  wire  m_394_io_x1; // @[MUL.scala 102:19]
  wire  m_394_io_x2; // @[MUL.scala 102:19]
  wire  m_394_io_x3; // @[MUL.scala 102:19]
  wire  m_394_io_s; // @[MUL.scala 102:19]
  wire  m_394_io_cout; // @[MUL.scala 102:19]
  wire  m_395_io_x1; // @[MUL.scala 102:19]
  wire  m_395_io_x2; // @[MUL.scala 102:19]
  wire  m_395_io_x3; // @[MUL.scala 102:19]
  wire  m_395_io_s; // @[MUL.scala 102:19]
  wire  m_395_io_cout; // @[MUL.scala 102:19]
  wire  m_396_io_x1; // @[MUL.scala 102:19]
  wire  m_396_io_x2; // @[MUL.scala 102:19]
  wire  m_396_io_x3; // @[MUL.scala 102:19]
  wire  m_396_io_s; // @[MUL.scala 102:19]
  wire  m_396_io_cout; // @[MUL.scala 102:19]
  wire  m_397_io_x1; // @[MUL.scala 102:19]
  wire  m_397_io_x2; // @[MUL.scala 102:19]
  wire  m_397_io_x3; // @[MUL.scala 102:19]
  wire  m_397_io_s; // @[MUL.scala 102:19]
  wire  m_397_io_cout; // @[MUL.scala 102:19]
  wire  m_398_io_x1; // @[MUL.scala 102:19]
  wire  m_398_io_x2; // @[MUL.scala 102:19]
  wire  m_398_io_x3; // @[MUL.scala 102:19]
  wire  m_398_io_s; // @[MUL.scala 102:19]
  wire  m_398_io_cout; // @[MUL.scala 102:19]
  wire  m_399_io_x1; // @[MUL.scala 102:19]
  wire  m_399_io_x2; // @[MUL.scala 102:19]
  wire  m_399_io_x3; // @[MUL.scala 102:19]
  wire  m_399_io_s; // @[MUL.scala 102:19]
  wire  m_399_io_cout; // @[MUL.scala 102:19]
  wire  m_400_io_x1; // @[MUL.scala 102:19]
  wire  m_400_io_x2; // @[MUL.scala 102:19]
  wire  m_400_io_x3; // @[MUL.scala 102:19]
  wire  m_400_io_s; // @[MUL.scala 102:19]
  wire  m_400_io_cout; // @[MUL.scala 102:19]
  wire  m_401_io_in_0; // @[MUL.scala 124:19]
  wire  m_401_io_in_1; // @[MUL.scala 124:19]
  wire  m_401_io_out_0; // @[MUL.scala 124:19]
  wire  m_401_io_out_1; // @[MUL.scala 124:19]
  wire  m_402_io_x1; // @[MUL.scala 102:19]
  wire  m_402_io_x2; // @[MUL.scala 102:19]
  wire  m_402_io_x3; // @[MUL.scala 102:19]
  wire  m_402_io_s; // @[MUL.scala 102:19]
  wire  m_402_io_cout; // @[MUL.scala 102:19]
  wire  m_403_io_in_0; // @[MUL.scala 124:19]
  wire  m_403_io_in_1; // @[MUL.scala 124:19]
  wire  m_403_io_out_0; // @[MUL.scala 124:19]
  wire  m_403_io_out_1; // @[MUL.scala 124:19]
  wire  m_404_io_x1; // @[MUL.scala 102:19]
  wire  m_404_io_x2; // @[MUL.scala 102:19]
  wire  m_404_io_x3; // @[MUL.scala 102:19]
  wire  m_404_io_s; // @[MUL.scala 102:19]
  wire  m_404_io_cout; // @[MUL.scala 102:19]
  wire  m_405_io_in_0; // @[MUL.scala 124:19]
  wire  m_405_io_in_1; // @[MUL.scala 124:19]
  wire  m_405_io_out_0; // @[MUL.scala 124:19]
  wire  m_405_io_out_1; // @[MUL.scala 124:19]
  wire  m_406_io_x1; // @[MUL.scala 102:19]
  wire  m_406_io_x2; // @[MUL.scala 102:19]
  wire  m_406_io_x3; // @[MUL.scala 102:19]
  wire  m_406_io_s; // @[MUL.scala 102:19]
  wire  m_406_io_cout; // @[MUL.scala 102:19]
  wire  m_407_io_in_0; // @[MUL.scala 124:19]
  wire  m_407_io_in_1; // @[MUL.scala 124:19]
  wire  m_407_io_out_0; // @[MUL.scala 124:19]
  wire  m_407_io_out_1; // @[MUL.scala 124:19]
  wire  m_408_io_x1; // @[MUL.scala 102:19]
  wire  m_408_io_x2; // @[MUL.scala 102:19]
  wire  m_408_io_x3; // @[MUL.scala 102:19]
  wire  m_408_io_s; // @[MUL.scala 102:19]
  wire  m_408_io_cout; // @[MUL.scala 102:19]
  wire  m_409_io_x1; // @[MUL.scala 102:19]
  wire  m_409_io_x2; // @[MUL.scala 102:19]
  wire  m_409_io_x3; // @[MUL.scala 102:19]
  wire  m_409_io_s; // @[MUL.scala 102:19]
  wire  m_409_io_cout; // @[MUL.scala 102:19]
  wire  m_410_io_x1; // @[MUL.scala 102:19]
  wire  m_410_io_x2; // @[MUL.scala 102:19]
  wire  m_410_io_x3; // @[MUL.scala 102:19]
  wire  m_410_io_s; // @[MUL.scala 102:19]
  wire  m_410_io_cout; // @[MUL.scala 102:19]
  wire  m_411_io_x1; // @[MUL.scala 102:19]
  wire  m_411_io_x2; // @[MUL.scala 102:19]
  wire  m_411_io_x3; // @[MUL.scala 102:19]
  wire  m_411_io_s; // @[MUL.scala 102:19]
  wire  m_411_io_cout; // @[MUL.scala 102:19]
  wire  m_412_io_x1; // @[MUL.scala 102:19]
  wire  m_412_io_x2; // @[MUL.scala 102:19]
  wire  m_412_io_x3; // @[MUL.scala 102:19]
  wire  m_412_io_s; // @[MUL.scala 102:19]
  wire  m_412_io_cout; // @[MUL.scala 102:19]
  wire  m_413_io_x1; // @[MUL.scala 102:19]
  wire  m_413_io_x2; // @[MUL.scala 102:19]
  wire  m_413_io_x3; // @[MUL.scala 102:19]
  wire  m_413_io_s; // @[MUL.scala 102:19]
  wire  m_413_io_cout; // @[MUL.scala 102:19]
  wire  m_414_io_x1; // @[MUL.scala 102:19]
  wire  m_414_io_x2; // @[MUL.scala 102:19]
  wire  m_414_io_x3; // @[MUL.scala 102:19]
  wire  m_414_io_s; // @[MUL.scala 102:19]
  wire  m_414_io_cout; // @[MUL.scala 102:19]
  wire  m_415_io_x1; // @[MUL.scala 102:19]
  wire  m_415_io_x2; // @[MUL.scala 102:19]
  wire  m_415_io_x3; // @[MUL.scala 102:19]
  wire  m_415_io_s; // @[MUL.scala 102:19]
  wire  m_415_io_cout; // @[MUL.scala 102:19]
  wire  m_416_io_x1; // @[MUL.scala 102:19]
  wire  m_416_io_x2; // @[MUL.scala 102:19]
  wire  m_416_io_x3; // @[MUL.scala 102:19]
  wire  m_416_io_s; // @[MUL.scala 102:19]
  wire  m_416_io_cout; // @[MUL.scala 102:19]
  wire  m_417_io_x1; // @[MUL.scala 102:19]
  wire  m_417_io_x2; // @[MUL.scala 102:19]
  wire  m_417_io_x3; // @[MUL.scala 102:19]
  wire  m_417_io_s; // @[MUL.scala 102:19]
  wire  m_417_io_cout; // @[MUL.scala 102:19]
  wire  m_418_io_x1; // @[MUL.scala 102:19]
  wire  m_418_io_x2; // @[MUL.scala 102:19]
  wire  m_418_io_x3; // @[MUL.scala 102:19]
  wire  m_418_io_s; // @[MUL.scala 102:19]
  wire  m_418_io_cout; // @[MUL.scala 102:19]
  wire  m_419_io_x1; // @[MUL.scala 102:19]
  wire  m_419_io_x2; // @[MUL.scala 102:19]
  wire  m_419_io_x3; // @[MUL.scala 102:19]
  wire  m_419_io_s; // @[MUL.scala 102:19]
  wire  m_419_io_cout; // @[MUL.scala 102:19]
  wire  m_420_io_x1; // @[MUL.scala 102:19]
  wire  m_420_io_x2; // @[MUL.scala 102:19]
  wire  m_420_io_x3; // @[MUL.scala 102:19]
  wire  m_420_io_s; // @[MUL.scala 102:19]
  wire  m_420_io_cout; // @[MUL.scala 102:19]
  wire  m_421_io_x1; // @[MUL.scala 102:19]
  wire  m_421_io_x2; // @[MUL.scala 102:19]
  wire  m_421_io_x3; // @[MUL.scala 102:19]
  wire  m_421_io_s; // @[MUL.scala 102:19]
  wire  m_421_io_cout; // @[MUL.scala 102:19]
  wire  m_422_io_x1; // @[MUL.scala 102:19]
  wire  m_422_io_x2; // @[MUL.scala 102:19]
  wire  m_422_io_x3; // @[MUL.scala 102:19]
  wire  m_422_io_s; // @[MUL.scala 102:19]
  wire  m_422_io_cout; // @[MUL.scala 102:19]
  wire  m_423_io_x1; // @[MUL.scala 102:19]
  wire  m_423_io_x2; // @[MUL.scala 102:19]
  wire  m_423_io_x3; // @[MUL.scala 102:19]
  wire  m_423_io_s; // @[MUL.scala 102:19]
  wire  m_423_io_cout; // @[MUL.scala 102:19]
  wire  m_424_io_x1; // @[MUL.scala 102:19]
  wire  m_424_io_x2; // @[MUL.scala 102:19]
  wire  m_424_io_x3; // @[MUL.scala 102:19]
  wire  m_424_io_s; // @[MUL.scala 102:19]
  wire  m_424_io_cout; // @[MUL.scala 102:19]
  wire  m_425_io_x1; // @[MUL.scala 102:19]
  wire  m_425_io_x2; // @[MUL.scala 102:19]
  wire  m_425_io_x3; // @[MUL.scala 102:19]
  wire  m_425_io_s; // @[MUL.scala 102:19]
  wire  m_425_io_cout; // @[MUL.scala 102:19]
  wire  m_426_io_x1; // @[MUL.scala 102:19]
  wire  m_426_io_x2; // @[MUL.scala 102:19]
  wire  m_426_io_x3; // @[MUL.scala 102:19]
  wire  m_426_io_s; // @[MUL.scala 102:19]
  wire  m_426_io_cout; // @[MUL.scala 102:19]
  wire  m_427_io_x1; // @[MUL.scala 102:19]
  wire  m_427_io_x2; // @[MUL.scala 102:19]
  wire  m_427_io_x3; // @[MUL.scala 102:19]
  wire  m_427_io_s; // @[MUL.scala 102:19]
  wire  m_427_io_cout; // @[MUL.scala 102:19]
  wire  m_428_io_in_0; // @[MUL.scala 124:19]
  wire  m_428_io_in_1; // @[MUL.scala 124:19]
  wire  m_428_io_out_0; // @[MUL.scala 124:19]
  wire  m_428_io_out_1; // @[MUL.scala 124:19]
  wire  m_429_io_x1; // @[MUL.scala 102:19]
  wire  m_429_io_x2; // @[MUL.scala 102:19]
  wire  m_429_io_x3; // @[MUL.scala 102:19]
  wire  m_429_io_s; // @[MUL.scala 102:19]
  wire  m_429_io_cout; // @[MUL.scala 102:19]
  wire  m_430_io_x1; // @[MUL.scala 102:19]
  wire  m_430_io_x2; // @[MUL.scala 102:19]
  wire  m_430_io_x3; // @[MUL.scala 102:19]
  wire  m_430_io_s; // @[MUL.scala 102:19]
  wire  m_430_io_cout; // @[MUL.scala 102:19]
  wire  m_431_io_in_0; // @[MUL.scala 124:19]
  wire  m_431_io_in_1; // @[MUL.scala 124:19]
  wire  m_431_io_out_0; // @[MUL.scala 124:19]
  wire  m_431_io_out_1; // @[MUL.scala 124:19]
  wire  m_432_io_x1; // @[MUL.scala 102:19]
  wire  m_432_io_x2; // @[MUL.scala 102:19]
  wire  m_432_io_x3; // @[MUL.scala 102:19]
  wire  m_432_io_s; // @[MUL.scala 102:19]
  wire  m_432_io_cout; // @[MUL.scala 102:19]
  wire  m_433_io_x1; // @[MUL.scala 102:19]
  wire  m_433_io_x2; // @[MUL.scala 102:19]
  wire  m_433_io_x3; // @[MUL.scala 102:19]
  wire  m_433_io_s; // @[MUL.scala 102:19]
  wire  m_433_io_cout; // @[MUL.scala 102:19]
  wire  m_434_io_in_0; // @[MUL.scala 124:19]
  wire  m_434_io_in_1; // @[MUL.scala 124:19]
  wire  m_434_io_out_0; // @[MUL.scala 124:19]
  wire  m_434_io_out_1; // @[MUL.scala 124:19]
  wire  m_435_io_x1; // @[MUL.scala 102:19]
  wire  m_435_io_x2; // @[MUL.scala 102:19]
  wire  m_435_io_x3; // @[MUL.scala 102:19]
  wire  m_435_io_s; // @[MUL.scala 102:19]
  wire  m_435_io_cout; // @[MUL.scala 102:19]
  wire  m_436_io_x1; // @[MUL.scala 102:19]
  wire  m_436_io_x2; // @[MUL.scala 102:19]
  wire  m_436_io_x3; // @[MUL.scala 102:19]
  wire  m_436_io_s; // @[MUL.scala 102:19]
  wire  m_436_io_cout; // @[MUL.scala 102:19]
  wire  m_437_io_in_0; // @[MUL.scala 124:19]
  wire  m_437_io_in_1; // @[MUL.scala 124:19]
  wire  m_437_io_out_0; // @[MUL.scala 124:19]
  wire  m_437_io_out_1; // @[MUL.scala 124:19]
  wire  m_438_io_x1; // @[MUL.scala 102:19]
  wire  m_438_io_x2; // @[MUL.scala 102:19]
  wire  m_438_io_x3; // @[MUL.scala 102:19]
  wire  m_438_io_s; // @[MUL.scala 102:19]
  wire  m_438_io_cout; // @[MUL.scala 102:19]
  wire  m_439_io_x1; // @[MUL.scala 102:19]
  wire  m_439_io_x2; // @[MUL.scala 102:19]
  wire  m_439_io_x3; // @[MUL.scala 102:19]
  wire  m_439_io_s; // @[MUL.scala 102:19]
  wire  m_439_io_cout; // @[MUL.scala 102:19]
  wire  m_440_io_in_0; // @[MUL.scala 124:19]
  wire  m_440_io_in_1; // @[MUL.scala 124:19]
  wire  m_440_io_out_0; // @[MUL.scala 124:19]
  wire  m_440_io_out_1; // @[MUL.scala 124:19]
  wire  m_441_io_x1; // @[MUL.scala 102:19]
  wire  m_441_io_x2; // @[MUL.scala 102:19]
  wire  m_441_io_x3; // @[MUL.scala 102:19]
  wire  m_441_io_s; // @[MUL.scala 102:19]
  wire  m_441_io_cout; // @[MUL.scala 102:19]
  wire  m_442_io_x1; // @[MUL.scala 102:19]
  wire  m_442_io_x2; // @[MUL.scala 102:19]
  wire  m_442_io_x3; // @[MUL.scala 102:19]
  wire  m_442_io_s; // @[MUL.scala 102:19]
  wire  m_442_io_cout; // @[MUL.scala 102:19]
  wire  m_443_io_in_0; // @[MUL.scala 124:19]
  wire  m_443_io_in_1; // @[MUL.scala 124:19]
  wire  m_443_io_out_0; // @[MUL.scala 124:19]
  wire  m_443_io_out_1; // @[MUL.scala 124:19]
  wire  m_444_io_x1; // @[MUL.scala 102:19]
  wire  m_444_io_x2; // @[MUL.scala 102:19]
  wire  m_444_io_x3; // @[MUL.scala 102:19]
  wire  m_444_io_s; // @[MUL.scala 102:19]
  wire  m_444_io_cout; // @[MUL.scala 102:19]
  wire  m_445_io_x1; // @[MUL.scala 102:19]
  wire  m_445_io_x2; // @[MUL.scala 102:19]
  wire  m_445_io_x3; // @[MUL.scala 102:19]
  wire  m_445_io_s; // @[MUL.scala 102:19]
  wire  m_445_io_cout; // @[MUL.scala 102:19]
  wire  m_446_io_in_0; // @[MUL.scala 124:19]
  wire  m_446_io_in_1; // @[MUL.scala 124:19]
  wire  m_446_io_out_0; // @[MUL.scala 124:19]
  wire  m_446_io_out_1; // @[MUL.scala 124:19]
  wire  m_447_io_x1; // @[MUL.scala 102:19]
  wire  m_447_io_x2; // @[MUL.scala 102:19]
  wire  m_447_io_x3; // @[MUL.scala 102:19]
  wire  m_447_io_s; // @[MUL.scala 102:19]
  wire  m_447_io_cout; // @[MUL.scala 102:19]
  wire  m_448_io_x1; // @[MUL.scala 102:19]
  wire  m_448_io_x2; // @[MUL.scala 102:19]
  wire  m_448_io_x3; // @[MUL.scala 102:19]
  wire  m_448_io_s; // @[MUL.scala 102:19]
  wire  m_448_io_cout; // @[MUL.scala 102:19]
  wire  m_449_io_in_0; // @[MUL.scala 124:19]
  wire  m_449_io_in_1; // @[MUL.scala 124:19]
  wire  m_449_io_out_0; // @[MUL.scala 124:19]
  wire  m_449_io_out_1; // @[MUL.scala 124:19]
  wire  m_450_io_x1; // @[MUL.scala 102:19]
  wire  m_450_io_x2; // @[MUL.scala 102:19]
  wire  m_450_io_x3; // @[MUL.scala 102:19]
  wire  m_450_io_s; // @[MUL.scala 102:19]
  wire  m_450_io_cout; // @[MUL.scala 102:19]
  wire  m_451_io_x1; // @[MUL.scala 102:19]
  wire  m_451_io_x2; // @[MUL.scala 102:19]
  wire  m_451_io_x3; // @[MUL.scala 102:19]
  wire  m_451_io_s; // @[MUL.scala 102:19]
  wire  m_451_io_cout; // @[MUL.scala 102:19]
  wire  m_452_io_in_0; // @[MUL.scala 124:19]
  wire  m_452_io_in_1; // @[MUL.scala 124:19]
  wire  m_452_io_out_0; // @[MUL.scala 124:19]
  wire  m_452_io_out_1; // @[MUL.scala 124:19]
  wire  m_453_io_x1; // @[MUL.scala 102:19]
  wire  m_453_io_x2; // @[MUL.scala 102:19]
  wire  m_453_io_x3; // @[MUL.scala 102:19]
  wire  m_453_io_s; // @[MUL.scala 102:19]
  wire  m_453_io_cout; // @[MUL.scala 102:19]
  wire  m_454_io_x1; // @[MUL.scala 102:19]
  wire  m_454_io_x2; // @[MUL.scala 102:19]
  wire  m_454_io_x3; // @[MUL.scala 102:19]
  wire  m_454_io_s; // @[MUL.scala 102:19]
  wire  m_454_io_cout; // @[MUL.scala 102:19]
  wire  m_455_io_in_0; // @[MUL.scala 124:19]
  wire  m_455_io_in_1; // @[MUL.scala 124:19]
  wire  m_455_io_out_0; // @[MUL.scala 124:19]
  wire  m_455_io_out_1; // @[MUL.scala 124:19]
  wire  m_456_io_x1; // @[MUL.scala 102:19]
  wire  m_456_io_x2; // @[MUL.scala 102:19]
  wire  m_456_io_x3; // @[MUL.scala 102:19]
  wire  m_456_io_s; // @[MUL.scala 102:19]
  wire  m_456_io_cout; // @[MUL.scala 102:19]
  wire  m_457_io_x1; // @[MUL.scala 102:19]
  wire  m_457_io_x2; // @[MUL.scala 102:19]
  wire  m_457_io_x3; // @[MUL.scala 102:19]
  wire  m_457_io_s; // @[MUL.scala 102:19]
  wire  m_457_io_cout; // @[MUL.scala 102:19]
  wire  m_458_io_x1; // @[MUL.scala 102:19]
  wire  m_458_io_x2; // @[MUL.scala 102:19]
  wire  m_458_io_x3; // @[MUL.scala 102:19]
  wire  m_458_io_s; // @[MUL.scala 102:19]
  wire  m_458_io_cout; // @[MUL.scala 102:19]
  wire  m_459_io_x1; // @[MUL.scala 102:19]
  wire  m_459_io_x2; // @[MUL.scala 102:19]
  wire  m_459_io_x3; // @[MUL.scala 102:19]
  wire  m_459_io_s; // @[MUL.scala 102:19]
  wire  m_459_io_cout; // @[MUL.scala 102:19]
  wire  m_460_io_x1; // @[MUL.scala 102:19]
  wire  m_460_io_x2; // @[MUL.scala 102:19]
  wire  m_460_io_x3; // @[MUL.scala 102:19]
  wire  m_460_io_s; // @[MUL.scala 102:19]
  wire  m_460_io_cout; // @[MUL.scala 102:19]
  wire  m_461_io_x1; // @[MUL.scala 102:19]
  wire  m_461_io_x2; // @[MUL.scala 102:19]
  wire  m_461_io_x3; // @[MUL.scala 102:19]
  wire  m_461_io_s; // @[MUL.scala 102:19]
  wire  m_461_io_cout; // @[MUL.scala 102:19]
  wire  m_462_io_x1; // @[MUL.scala 102:19]
  wire  m_462_io_x2; // @[MUL.scala 102:19]
  wire  m_462_io_x3; // @[MUL.scala 102:19]
  wire  m_462_io_s; // @[MUL.scala 102:19]
  wire  m_462_io_cout; // @[MUL.scala 102:19]
  wire  m_463_io_x1; // @[MUL.scala 102:19]
  wire  m_463_io_x2; // @[MUL.scala 102:19]
  wire  m_463_io_x3; // @[MUL.scala 102:19]
  wire  m_463_io_s; // @[MUL.scala 102:19]
  wire  m_463_io_cout; // @[MUL.scala 102:19]
  wire  m_464_io_x1; // @[MUL.scala 102:19]
  wire  m_464_io_x2; // @[MUL.scala 102:19]
  wire  m_464_io_x3; // @[MUL.scala 102:19]
  wire  m_464_io_s; // @[MUL.scala 102:19]
  wire  m_464_io_cout; // @[MUL.scala 102:19]
  wire  m_465_io_x1; // @[MUL.scala 102:19]
  wire  m_465_io_x2; // @[MUL.scala 102:19]
  wire  m_465_io_x3; // @[MUL.scala 102:19]
  wire  m_465_io_s; // @[MUL.scala 102:19]
  wire  m_465_io_cout; // @[MUL.scala 102:19]
  wire  m_466_io_x1; // @[MUL.scala 102:19]
  wire  m_466_io_x2; // @[MUL.scala 102:19]
  wire  m_466_io_x3; // @[MUL.scala 102:19]
  wire  m_466_io_s; // @[MUL.scala 102:19]
  wire  m_466_io_cout; // @[MUL.scala 102:19]
  wire  m_467_io_x1; // @[MUL.scala 102:19]
  wire  m_467_io_x2; // @[MUL.scala 102:19]
  wire  m_467_io_x3; // @[MUL.scala 102:19]
  wire  m_467_io_s; // @[MUL.scala 102:19]
  wire  m_467_io_cout; // @[MUL.scala 102:19]
  wire  m_468_io_x1; // @[MUL.scala 102:19]
  wire  m_468_io_x2; // @[MUL.scala 102:19]
  wire  m_468_io_x3; // @[MUL.scala 102:19]
  wire  m_468_io_s; // @[MUL.scala 102:19]
  wire  m_468_io_cout; // @[MUL.scala 102:19]
  wire  m_469_io_x1; // @[MUL.scala 102:19]
  wire  m_469_io_x2; // @[MUL.scala 102:19]
  wire  m_469_io_x3; // @[MUL.scala 102:19]
  wire  m_469_io_s; // @[MUL.scala 102:19]
  wire  m_469_io_cout; // @[MUL.scala 102:19]
  wire  m_470_io_x1; // @[MUL.scala 102:19]
  wire  m_470_io_x2; // @[MUL.scala 102:19]
  wire  m_470_io_x3; // @[MUL.scala 102:19]
  wire  m_470_io_s; // @[MUL.scala 102:19]
  wire  m_470_io_cout; // @[MUL.scala 102:19]
  wire  m_471_io_x1; // @[MUL.scala 102:19]
  wire  m_471_io_x2; // @[MUL.scala 102:19]
  wire  m_471_io_x3; // @[MUL.scala 102:19]
  wire  m_471_io_s; // @[MUL.scala 102:19]
  wire  m_471_io_cout; // @[MUL.scala 102:19]
  wire  m_472_io_x1; // @[MUL.scala 102:19]
  wire  m_472_io_x2; // @[MUL.scala 102:19]
  wire  m_472_io_x3; // @[MUL.scala 102:19]
  wire  m_472_io_s; // @[MUL.scala 102:19]
  wire  m_472_io_cout; // @[MUL.scala 102:19]
  wire  m_473_io_x1; // @[MUL.scala 102:19]
  wire  m_473_io_x2; // @[MUL.scala 102:19]
  wire  m_473_io_x3; // @[MUL.scala 102:19]
  wire  m_473_io_s; // @[MUL.scala 102:19]
  wire  m_473_io_cout; // @[MUL.scala 102:19]
  wire  m_474_io_x1; // @[MUL.scala 102:19]
  wire  m_474_io_x2; // @[MUL.scala 102:19]
  wire  m_474_io_x3; // @[MUL.scala 102:19]
  wire  m_474_io_s; // @[MUL.scala 102:19]
  wire  m_474_io_cout; // @[MUL.scala 102:19]
  wire  m_475_io_x1; // @[MUL.scala 102:19]
  wire  m_475_io_x2; // @[MUL.scala 102:19]
  wire  m_475_io_x3; // @[MUL.scala 102:19]
  wire  m_475_io_s; // @[MUL.scala 102:19]
  wire  m_475_io_cout; // @[MUL.scala 102:19]
  wire  m_476_io_x1; // @[MUL.scala 102:19]
  wire  m_476_io_x2; // @[MUL.scala 102:19]
  wire  m_476_io_x3; // @[MUL.scala 102:19]
  wire  m_476_io_s; // @[MUL.scala 102:19]
  wire  m_476_io_cout; // @[MUL.scala 102:19]
  wire  m_477_io_x1; // @[MUL.scala 102:19]
  wire  m_477_io_x2; // @[MUL.scala 102:19]
  wire  m_477_io_x3; // @[MUL.scala 102:19]
  wire  m_477_io_s; // @[MUL.scala 102:19]
  wire  m_477_io_cout; // @[MUL.scala 102:19]
  wire  m_478_io_x1; // @[MUL.scala 102:19]
  wire  m_478_io_x2; // @[MUL.scala 102:19]
  wire  m_478_io_x3; // @[MUL.scala 102:19]
  wire  m_478_io_s; // @[MUL.scala 102:19]
  wire  m_478_io_cout; // @[MUL.scala 102:19]
  wire  m_479_io_x1; // @[MUL.scala 102:19]
  wire  m_479_io_x2; // @[MUL.scala 102:19]
  wire  m_479_io_x3; // @[MUL.scala 102:19]
  wire  m_479_io_s; // @[MUL.scala 102:19]
  wire  m_479_io_cout; // @[MUL.scala 102:19]
  wire  m_480_io_x1; // @[MUL.scala 102:19]
  wire  m_480_io_x2; // @[MUL.scala 102:19]
  wire  m_480_io_x3; // @[MUL.scala 102:19]
  wire  m_480_io_s; // @[MUL.scala 102:19]
  wire  m_480_io_cout; // @[MUL.scala 102:19]
  wire  m_481_io_x1; // @[MUL.scala 102:19]
  wire  m_481_io_x2; // @[MUL.scala 102:19]
  wire  m_481_io_x3; // @[MUL.scala 102:19]
  wire  m_481_io_s; // @[MUL.scala 102:19]
  wire  m_481_io_cout; // @[MUL.scala 102:19]
  wire  m_482_io_x1; // @[MUL.scala 102:19]
  wire  m_482_io_x2; // @[MUL.scala 102:19]
  wire  m_482_io_x3; // @[MUL.scala 102:19]
  wire  m_482_io_s; // @[MUL.scala 102:19]
  wire  m_482_io_cout; // @[MUL.scala 102:19]
  wire  m_483_io_x1; // @[MUL.scala 102:19]
  wire  m_483_io_x2; // @[MUL.scala 102:19]
  wire  m_483_io_x3; // @[MUL.scala 102:19]
  wire  m_483_io_s; // @[MUL.scala 102:19]
  wire  m_483_io_cout; // @[MUL.scala 102:19]
  wire  m_484_io_x1; // @[MUL.scala 102:19]
  wire  m_484_io_x2; // @[MUL.scala 102:19]
  wire  m_484_io_x3; // @[MUL.scala 102:19]
  wire  m_484_io_s; // @[MUL.scala 102:19]
  wire  m_484_io_cout; // @[MUL.scala 102:19]
  wire  m_485_io_x1; // @[MUL.scala 102:19]
  wire  m_485_io_x2; // @[MUL.scala 102:19]
  wire  m_485_io_x3; // @[MUL.scala 102:19]
  wire  m_485_io_s; // @[MUL.scala 102:19]
  wire  m_485_io_cout; // @[MUL.scala 102:19]
  wire  m_486_io_x1; // @[MUL.scala 102:19]
  wire  m_486_io_x2; // @[MUL.scala 102:19]
  wire  m_486_io_x3; // @[MUL.scala 102:19]
  wire  m_486_io_s; // @[MUL.scala 102:19]
  wire  m_486_io_cout; // @[MUL.scala 102:19]
  wire  m_487_io_x1; // @[MUL.scala 102:19]
  wire  m_487_io_x2; // @[MUL.scala 102:19]
  wire  m_487_io_x3; // @[MUL.scala 102:19]
  wire  m_487_io_s; // @[MUL.scala 102:19]
  wire  m_487_io_cout; // @[MUL.scala 102:19]
  wire  m_488_io_x1; // @[MUL.scala 102:19]
  wire  m_488_io_x2; // @[MUL.scala 102:19]
  wire  m_488_io_x3; // @[MUL.scala 102:19]
  wire  m_488_io_s; // @[MUL.scala 102:19]
  wire  m_488_io_cout; // @[MUL.scala 102:19]
  wire  m_489_io_in_0; // @[MUL.scala 124:19]
  wire  m_489_io_in_1; // @[MUL.scala 124:19]
  wire  m_489_io_out_0; // @[MUL.scala 124:19]
  wire  m_489_io_out_1; // @[MUL.scala 124:19]
  wire  m_490_io_in_0; // @[MUL.scala 124:19]
  wire  m_490_io_in_1; // @[MUL.scala 124:19]
  wire  m_490_io_out_0; // @[MUL.scala 124:19]
  wire  m_490_io_out_1; // @[MUL.scala 124:19]
  wire  m_491_io_in_0; // @[MUL.scala 124:19]
  wire  m_491_io_in_1; // @[MUL.scala 124:19]
  wire  m_491_io_out_0; // @[MUL.scala 124:19]
  wire  m_491_io_out_1; // @[MUL.scala 124:19]
  wire  m_492_io_in_0; // @[MUL.scala 124:19]
  wire  m_492_io_in_1; // @[MUL.scala 124:19]
  wire  m_492_io_out_0; // @[MUL.scala 124:19]
  wire  m_492_io_out_1; // @[MUL.scala 124:19]
  wire  m_493_io_in_0; // @[MUL.scala 124:19]
  wire  m_493_io_in_1; // @[MUL.scala 124:19]
  wire  m_493_io_out_0; // @[MUL.scala 124:19]
  wire  m_493_io_out_1; // @[MUL.scala 124:19]
  wire  m_494_io_in_0; // @[MUL.scala 124:19]
  wire  m_494_io_in_1; // @[MUL.scala 124:19]
  wire  m_494_io_out_0; // @[MUL.scala 124:19]
  wire  m_494_io_out_1; // @[MUL.scala 124:19]
  wire  m_495_io_in_0; // @[MUL.scala 124:19]
  wire  m_495_io_in_1; // @[MUL.scala 124:19]
  wire  m_495_io_out_0; // @[MUL.scala 124:19]
  wire  m_495_io_out_1; // @[MUL.scala 124:19]
  wire  m_496_io_in_0; // @[MUL.scala 124:19]
  wire  m_496_io_in_1; // @[MUL.scala 124:19]
  wire  m_496_io_out_0; // @[MUL.scala 124:19]
  wire  m_496_io_out_1; // @[MUL.scala 124:19]
  wire  m_497_io_in_0; // @[MUL.scala 124:19]
  wire  m_497_io_in_1; // @[MUL.scala 124:19]
  wire  m_497_io_out_0; // @[MUL.scala 124:19]
  wire  m_497_io_out_1; // @[MUL.scala 124:19]
  wire  m_498_io_in_0; // @[MUL.scala 124:19]
  wire  m_498_io_in_1; // @[MUL.scala 124:19]
  wire  m_498_io_out_0; // @[MUL.scala 124:19]
  wire  m_498_io_out_1; // @[MUL.scala 124:19]
  wire  m_499_io_in_0; // @[MUL.scala 124:19]
  wire  m_499_io_in_1; // @[MUL.scala 124:19]
  wire  m_499_io_out_0; // @[MUL.scala 124:19]
  wire  m_499_io_out_1; // @[MUL.scala 124:19]
  wire  m_500_io_in_0; // @[MUL.scala 124:19]
  wire  m_500_io_in_1; // @[MUL.scala 124:19]
  wire  m_500_io_out_0; // @[MUL.scala 124:19]
  wire  m_500_io_out_1; // @[MUL.scala 124:19]
  wire  m_501_io_in_0; // @[MUL.scala 124:19]
  wire  m_501_io_in_1; // @[MUL.scala 124:19]
  wire  m_501_io_out_0; // @[MUL.scala 124:19]
  wire  m_501_io_out_1; // @[MUL.scala 124:19]
  wire  m_502_io_in_0; // @[MUL.scala 124:19]
  wire  m_502_io_in_1; // @[MUL.scala 124:19]
  wire  m_502_io_out_0; // @[MUL.scala 124:19]
  wire  m_502_io_out_1; // @[MUL.scala 124:19]
  wire  m_503_io_x1; // @[MUL.scala 102:19]
  wire  m_503_io_x2; // @[MUL.scala 102:19]
  wire  m_503_io_x3; // @[MUL.scala 102:19]
  wire  m_503_io_s; // @[MUL.scala 102:19]
  wire  m_503_io_cout; // @[MUL.scala 102:19]
  wire  m_504_io_x1; // @[MUL.scala 102:19]
  wire  m_504_io_x2; // @[MUL.scala 102:19]
  wire  m_504_io_x3; // @[MUL.scala 102:19]
  wire  m_504_io_s; // @[MUL.scala 102:19]
  wire  m_504_io_cout; // @[MUL.scala 102:19]
  wire  m_505_io_x1; // @[MUL.scala 102:19]
  wire  m_505_io_x2; // @[MUL.scala 102:19]
  wire  m_505_io_x3; // @[MUL.scala 102:19]
  wire  m_505_io_s; // @[MUL.scala 102:19]
  wire  m_505_io_cout; // @[MUL.scala 102:19]
  wire  m_506_io_x1; // @[MUL.scala 102:19]
  wire  m_506_io_x2; // @[MUL.scala 102:19]
  wire  m_506_io_x3; // @[MUL.scala 102:19]
  wire  m_506_io_s; // @[MUL.scala 102:19]
  wire  m_506_io_cout; // @[MUL.scala 102:19]
  wire  m_507_io_x1; // @[MUL.scala 102:19]
  wire  m_507_io_x2; // @[MUL.scala 102:19]
  wire  m_507_io_x3; // @[MUL.scala 102:19]
  wire  m_507_io_s; // @[MUL.scala 102:19]
  wire  m_507_io_cout; // @[MUL.scala 102:19]
  wire  m_508_io_x1; // @[MUL.scala 102:19]
  wire  m_508_io_x2; // @[MUL.scala 102:19]
  wire  m_508_io_x3; // @[MUL.scala 102:19]
  wire  m_508_io_s; // @[MUL.scala 102:19]
  wire  m_508_io_cout; // @[MUL.scala 102:19]
  wire  m_509_io_x1; // @[MUL.scala 102:19]
  wire  m_509_io_x2; // @[MUL.scala 102:19]
  wire  m_509_io_x3; // @[MUL.scala 102:19]
  wire  m_509_io_s; // @[MUL.scala 102:19]
  wire  m_509_io_cout; // @[MUL.scala 102:19]
  wire  m_510_io_x1; // @[MUL.scala 102:19]
  wire  m_510_io_x2; // @[MUL.scala 102:19]
  wire  m_510_io_x3; // @[MUL.scala 102:19]
  wire  m_510_io_s; // @[MUL.scala 102:19]
  wire  m_510_io_cout; // @[MUL.scala 102:19]
  wire  m_511_io_x1; // @[MUL.scala 102:19]
  wire  m_511_io_x2; // @[MUL.scala 102:19]
  wire  m_511_io_x3; // @[MUL.scala 102:19]
  wire  m_511_io_s; // @[MUL.scala 102:19]
  wire  m_511_io_cout; // @[MUL.scala 102:19]
  wire  m_512_io_x1; // @[MUL.scala 102:19]
  wire  m_512_io_x2; // @[MUL.scala 102:19]
  wire  m_512_io_x3; // @[MUL.scala 102:19]
  wire  m_512_io_s; // @[MUL.scala 102:19]
  wire  m_512_io_cout; // @[MUL.scala 102:19]
  wire  m_513_io_x1; // @[MUL.scala 102:19]
  wire  m_513_io_x2; // @[MUL.scala 102:19]
  wire  m_513_io_x3; // @[MUL.scala 102:19]
  wire  m_513_io_s; // @[MUL.scala 102:19]
  wire  m_513_io_cout; // @[MUL.scala 102:19]
  wire  m_514_io_x1; // @[MUL.scala 102:19]
  wire  m_514_io_x2; // @[MUL.scala 102:19]
  wire  m_514_io_x3; // @[MUL.scala 102:19]
  wire  m_514_io_s; // @[MUL.scala 102:19]
  wire  m_514_io_cout; // @[MUL.scala 102:19]
  wire  m_515_io_x1; // @[MUL.scala 102:19]
  wire  m_515_io_x2; // @[MUL.scala 102:19]
  wire  m_515_io_x3; // @[MUL.scala 102:19]
  wire  m_515_io_s; // @[MUL.scala 102:19]
  wire  m_515_io_cout; // @[MUL.scala 102:19]
  wire  m_516_io_x1; // @[MUL.scala 102:19]
  wire  m_516_io_x2; // @[MUL.scala 102:19]
  wire  m_516_io_x3; // @[MUL.scala 102:19]
  wire  m_516_io_s; // @[MUL.scala 102:19]
  wire  m_516_io_cout; // @[MUL.scala 102:19]
  wire  m_517_io_x1; // @[MUL.scala 102:19]
  wire  m_517_io_x2; // @[MUL.scala 102:19]
  wire  m_517_io_x3; // @[MUL.scala 102:19]
  wire  m_517_io_s; // @[MUL.scala 102:19]
  wire  m_517_io_cout; // @[MUL.scala 102:19]
  wire  m_518_io_in_0; // @[MUL.scala 124:19]
  wire  m_518_io_in_1; // @[MUL.scala 124:19]
  wire  m_518_io_out_0; // @[MUL.scala 124:19]
  wire  m_518_io_out_1; // @[MUL.scala 124:19]
  wire  m_519_io_x1; // @[MUL.scala 102:19]
  wire  m_519_io_x2; // @[MUL.scala 102:19]
  wire  m_519_io_x3; // @[MUL.scala 102:19]
  wire  m_519_io_s; // @[MUL.scala 102:19]
  wire  m_519_io_cout; // @[MUL.scala 102:19]
  wire  m_520_io_in_0; // @[MUL.scala 124:19]
  wire  m_520_io_in_1; // @[MUL.scala 124:19]
  wire  m_520_io_out_0; // @[MUL.scala 124:19]
  wire  m_520_io_out_1; // @[MUL.scala 124:19]
  wire  m_521_io_x1; // @[MUL.scala 102:19]
  wire  m_521_io_x2; // @[MUL.scala 102:19]
  wire  m_521_io_x3; // @[MUL.scala 102:19]
  wire  m_521_io_s; // @[MUL.scala 102:19]
  wire  m_521_io_cout; // @[MUL.scala 102:19]
  wire  m_522_io_in_0; // @[MUL.scala 124:19]
  wire  m_522_io_in_1; // @[MUL.scala 124:19]
  wire  m_522_io_out_0; // @[MUL.scala 124:19]
  wire  m_522_io_out_1; // @[MUL.scala 124:19]
  wire  m_523_io_x1; // @[MUL.scala 102:19]
  wire  m_523_io_x2; // @[MUL.scala 102:19]
  wire  m_523_io_x3; // @[MUL.scala 102:19]
  wire  m_523_io_s; // @[MUL.scala 102:19]
  wire  m_523_io_cout; // @[MUL.scala 102:19]
  wire  m_524_io_in_0; // @[MUL.scala 124:19]
  wire  m_524_io_in_1; // @[MUL.scala 124:19]
  wire  m_524_io_out_0; // @[MUL.scala 124:19]
  wire  m_524_io_out_1; // @[MUL.scala 124:19]
  wire  m_525_io_x1; // @[MUL.scala 102:19]
  wire  m_525_io_x2; // @[MUL.scala 102:19]
  wire  m_525_io_x3; // @[MUL.scala 102:19]
  wire  m_525_io_s; // @[MUL.scala 102:19]
  wire  m_525_io_cout; // @[MUL.scala 102:19]
  wire  m_526_io_in_0; // @[MUL.scala 124:19]
  wire  m_526_io_in_1; // @[MUL.scala 124:19]
  wire  m_526_io_out_0; // @[MUL.scala 124:19]
  wire  m_526_io_out_1; // @[MUL.scala 124:19]
  wire  m_527_io_x1; // @[MUL.scala 102:19]
  wire  m_527_io_x2; // @[MUL.scala 102:19]
  wire  m_527_io_x3; // @[MUL.scala 102:19]
  wire  m_527_io_s; // @[MUL.scala 102:19]
  wire  m_527_io_cout; // @[MUL.scala 102:19]
  wire  m_528_io_x1; // @[MUL.scala 102:19]
  wire  m_528_io_x2; // @[MUL.scala 102:19]
  wire  m_528_io_x3; // @[MUL.scala 102:19]
  wire  m_528_io_s; // @[MUL.scala 102:19]
  wire  m_528_io_cout; // @[MUL.scala 102:19]
  wire  m_529_io_x1; // @[MUL.scala 102:19]
  wire  m_529_io_x2; // @[MUL.scala 102:19]
  wire  m_529_io_x3; // @[MUL.scala 102:19]
  wire  m_529_io_s; // @[MUL.scala 102:19]
  wire  m_529_io_cout; // @[MUL.scala 102:19]
  wire  m_530_io_x1; // @[MUL.scala 102:19]
  wire  m_530_io_x2; // @[MUL.scala 102:19]
  wire  m_530_io_x3; // @[MUL.scala 102:19]
  wire  m_530_io_s; // @[MUL.scala 102:19]
  wire  m_530_io_cout; // @[MUL.scala 102:19]
  wire  m_531_io_x1; // @[MUL.scala 102:19]
  wire  m_531_io_x2; // @[MUL.scala 102:19]
  wire  m_531_io_x3; // @[MUL.scala 102:19]
  wire  m_531_io_s; // @[MUL.scala 102:19]
  wire  m_531_io_cout; // @[MUL.scala 102:19]
  wire  m_532_io_x1; // @[MUL.scala 102:19]
  wire  m_532_io_x2; // @[MUL.scala 102:19]
  wire  m_532_io_x3; // @[MUL.scala 102:19]
  wire  m_532_io_s; // @[MUL.scala 102:19]
  wire  m_532_io_cout; // @[MUL.scala 102:19]
  wire  m_533_io_x1; // @[MUL.scala 102:19]
  wire  m_533_io_x2; // @[MUL.scala 102:19]
  wire  m_533_io_x3; // @[MUL.scala 102:19]
  wire  m_533_io_s; // @[MUL.scala 102:19]
  wire  m_533_io_cout; // @[MUL.scala 102:19]
  wire  m_534_io_x1; // @[MUL.scala 102:19]
  wire  m_534_io_x2; // @[MUL.scala 102:19]
  wire  m_534_io_x3; // @[MUL.scala 102:19]
  wire  m_534_io_s; // @[MUL.scala 102:19]
  wire  m_534_io_cout; // @[MUL.scala 102:19]
  wire  m_535_io_x1; // @[MUL.scala 102:19]
  wire  m_535_io_x2; // @[MUL.scala 102:19]
  wire  m_535_io_x3; // @[MUL.scala 102:19]
  wire  m_535_io_s; // @[MUL.scala 102:19]
  wire  m_535_io_cout; // @[MUL.scala 102:19]
  wire  m_536_io_x1; // @[MUL.scala 102:19]
  wire  m_536_io_x2; // @[MUL.scala 102:19]
  wire  m_536_io_x3; // @[MUL.scala 102:19]
  wire  m_536_io_s; // @[MUL.scala 102:19]
  wire  m_536_io_cout; // @[MUL.scala 102:19]
  wire  m_537_io_x1; // @[MUL.scala 102:19]
  wire  m_537_io_x2; // @[MUL.scala 102:19]
  wire  m_537_io_x3; // @[MUL.scala 102:19]
  wire  m_537_io_s; // @[MUL.scala 102:19]
  wire  m_537_io_cout; // @[MUL.scala 102:19]
  wire  m_538_io_x1; // @[MUL.scala 102:19]
  wire  m_538_io_x2; // @[MUL.scala 102:19]
  wire  m_538_io_x3; // @[MUL.scala 102:19]
  wire  m_538_io_s; // @[MUL.scala 102:19]
  wire  m_538_io_cout; // @[MUL.scala 102:19]
  wire  m_539_io_x1; // @[MUL.scala 102:19]
  wire  m_539_io_x2; // @[MUL.scala 102:19]
  wire  m_539_io_x3; // @[MUL.scala 102:19]
  wire  m_539_io_s; // @[MUL.scala 102:19]
  wire  m_539_io_cout; // @[MUL.scala 102:19]
  wire  m_540_io_x1; // @[MUL.scala 102:19]
  wire  m_540_io_x2; // @[MUL.scala 102:19]
  wire  m_540_io_x3; // @[MUL.scala 102:19]
  wire  m_540_io_s; // @[MUL.scala 102:19]
  wire  m_540_io_cout; // @[MUL.scala 102:19]
  wire  m_541_io_x1; // @[MUL.scala 102:19]
  wire  m_541_io_x2; // @[MUL.scala 102:19]
  wire  m_541_io_x3; // @[MUL.scala 102:19]
  wire  m_541_io_s; // @[MUL.scala 102:19]
  wire  m_541_io_cout; // @[MUL.scala 102:19]
  wire  m_542_io_x1; // @[MUL.scala 102:19]
  wire  m_542_io_x2; // @[MUL.scala 102:19]
  wire  m_542_io_x3; // @[MUL.scala 102:19]
  wire  m_542_io_s; // @[MUL.scala 102:19]
  wire  m_542_io_cout; // @[MUL.scala 102:19]
  wire  m_543_io_x1; // @[MUL.scala 102:19]
  wire  m_543_io_x2; // @[MUL.scala 102:19]
  wire  m_543_io_x3; // @[MUL.scala 102:19]
  wire  m_543_io_s; // @[MUL.scala 102:19]
  wire  m_543_io_cout; // @[MUL.scala 102:19]
  wire  m_544_io_x1; // @[MUL.scala 102:19]
  wire  m_544_io_x2; // @[MUL.scala 102:19]
  wire  m_544_io_x3; // @[MUL.scala 102:19]
  wire  m_544_io_s; // @[MUL.scala 102:19]
  wire  m_544_io_cout; // @[MUL.scala 102:19]
  wire  m_545_io_x1; // @[MUL.scala 102:19]
  wire  m_545_io_x2; // @[MUL.scala 102:19]
  wire  m_545_io_x3; // @[MUL.scala 102:19]
  wire  m_545_io_s; // @[MUL.scala 102:19]
  wire  m_545_io_cout; // @[MUL.scala 102:19]
  wire  m_546_io_x1; // @[MUL.scala 102:19]
  wire  m_546_io_x2; // @[MUL.scala 102:19]
  wire  m_546_io_x3; // @[MUL.scala 102:19]
  wire  m_546_io_s; // @[MUL.scala 102:19]
  wire  m_546_io_cout; // @[MUL.scala 102:19]
  wire  m_547_io_x1; // @[MUL.scala 102:19]
  wire  m_547_io_x2; // @[MUL.scala 102:19]
  wire  m_547_io_x3; // @[MUL.scala 102:19]
  wire  m_547_io_s; // @[MUL.scala 102:19]
  wire  m_547_io_cout; // @[MUL.scala 102:19]
  wire  m_548_io_in_0; // @[MUL.scala 124:19]
  wire  m_548_io_in_1; // @[MUL.scala 124:19]
  wire  m_548_io_out_0; // @[MUL.scala 124:19]
  wire  m_548_io_out_1; // @[MUL.scala 124:19]
  wire  m_549_io_x1; // @[MUL.scala 102:19]
  wire  m_549_io_x2; // @[MUL.scala 102:19]
  wire  m_549_io_x3; // @[MUL.scala 102:19]
  wire  m_549_io_s; // @[MUL.scala 102:19]
  wire  m_549_io_cout; // @[MUL.scala 102:19]
  wire  m_550_io_in_0; // @[MUL.scala 124:19]
  wire  m_550_io_in_1; // @[MUL.scala 124:19]
  wire  m_550_io_out_0; // @[MUL.scala 124:19]
  wire  m_550_io_out_1; // @[MUL.scala 124:19]
  wire  m_551_io_x1; // @[MUL.scala 102:19]
  wire  m_551_io_x2; // @[MUL.scala 102:19]
  wire  m_551_io_x3; // @[MUL.scala 102:19]
  wire  m_551_io_s; // @[MUL.scala 102:19]
  wire  m_551_io_cout; // @[MUL.scala 102:19]
  wire  m_552_io_in_0; // @[MUL.scala 124:19]
  wire  m_552_io_in_1; // @[MUL.scala 124:19]
  wire  m_552_io_out_0; // @[MUL.scala 124:19]
  wire  m_552_io_out_1; // @[MUL.scala 124:19]
  wire  m_553_io_x1; // @[MUL.scala 102:19]
  wire  m_553_io_x2; // @[MUL.scala 102:19]
  wire  m_553_io_x3; // @[MUL.scala 102:19]
  wire  m_553_io_s; // @[MUL.scala 102:19]
  wire  m_553_io_cout; // @[MUL.scala 102:19]
  wire  m_554_io_x1; // @[MUL.scala 102:19]
  wire  m_554_io_x2; // @[MUL.scala 102:19]
  wire  m_554_io_x3; // @[MUL.scala 102:19]
  wire  m_554_io_s; // @[MUL.scala 102:19]
  wire  m_554_io_cout; // @[MUL.scala 102:19]
  wire  m_555_io_x1; // @[MUL.scala 102:19]
  wire  m_555_io_x2; // @[MUL.scala 102:19]
  wire  m_555_io_x3; // @[MUL.scala 102:19]
  wire  m_555_io_s; // @[MUL.scala 102:19]
  wire  m_555_io_cout; // @[MUL.scala 102:19]
  wire  m_556_io_x1; // @[MUL.scala 102:19]
  wire  m_556_io_x2; // @[MUL.scala 102:19]
  wire  m_556_io_x3; // @[MUL.scala 102:19]
  wire  m_556_io_s; // @[MUL.scala 102:19]
  wire  m_556_io_cout; // @[MUL.scala 102:19]
  wire  m_557_io_x1; // @[MUL.scala 102:19]
  wire  m_557_io_x2; // @[MUL.scala 102:19]
  wire  m_557_io_x3; // @[MUL.scala 102:19]
  wire  m_557_io_s; // @[MUL.scala 102:19]
  wire  m_557_io_cout; // @[MUL.scala 102:19]
  wire  m_558_io_x1; // @[MUL.scala 102:19]
  wire  m_558_io_x2; // @[MUL.scala 102:19]
  wire  m_558_io_x3; // @[MUL.scala 102:19]
  wire  m_558_io_s; // @[MUL.scala 102:19]
  wire  m_558_io_cout; // @[MUL.scala 102:19]
  wire  m_559_io_x1; // @[MUL.scala 102:19]
  wire  m_559_io_x2; // @[MUL.scala 102:19]
  wire  m_559_io_x3; // @[MUL.scala 102:19]
  wire  m_559_io_s; // @[MUL.scala 102:19]
  wire  m_559_io_cout; // @[MUL.scala 102:19]
  wire  m_560_io_x1; // @[MUL.scala 102:19]
  wire  m_560_io_x2; // @[MUL.scala 102:19]
  wire  m_560_io_x3; // @[MUL.scala 102:19]
  wire  m_560_io_s; // @[MUL.scala 102:19]
  wire  m_560_io_cout; // @[MUL.scala 102:19]
  wire  m_561_io_x1; // @[MUL.scala 102:19]
  wire  m_561_io_x2; // @[MUL.scala 102:19]
  wire  m_561_io_x3; // @[MUL.scala 102:19]
  wire  m_561_io_s; // @[MUL.scala 102:19]
  wire  m_561_io_cout; // @[MUL.scala 102:19]
  wire  m_562_io_x1; // @[MUL.scala 102:19]
  wire  m_562_io_x2; // @[MUL.scala 102:19]
  wire  m_562_io_x3; // @[MUL.scala 102:19]
  wire  m_562_io_s; // @[MUL.scala 102:19]
  wire  m_562_io_cout; // @[MUL.scala 102:19]
  wire  m_563_io_x1; // @[MUL.scala 102:19]
  wire  m_563_io_x2; // @[MUL.scala 102:19]
  wire  m_563_io_x3; // @[MUL.scala 102:19]
  wire  m_563_io_s; // @[MUL.scala 102:19]
  wire  m_563_io_cout; // @[MUL.scala 102:19]
  wire  m_564_io_x1; // @[MUL.scala 102:19]
  wire  m_564_io_x2; // @[MUL.scala 102:19]
  wire  m_564_io_x3; // @[MUL.scala 102:19]
  wire  m_564_io_s; // @[MUL.scala 102:19]
  wire  m_564_io_cout; // @[MUL.scala 102:19]
  wire  m_565_io_x1; // @[MUL.scala 102:19]
  wire  m_565_io_x2; // @[MUL.scala 102:19]
  wire  m_565_io_x3; // @[MUL.scala 102:19]
  wire  m_565_io_s; // @[MUL.scala 102:19]
  wire  m_565_io_cout; // @[MUL.scala 102:19]
  wire  m_566_io_x1; // @[MUL.scala 102:19]
  wire  m_566_io_x2; // @[MUL.scala 102:19]
  wire  m_566_io_x3; // @[MUL.scala 102:19]
  wire  m_566_io_s; // @[MUL.scala 102:19]
  wire  m_566_io_cout; // @[MUL.scala 102:19]
  wire  m_567_io_in_0; // @[MUL.scala 124:19]
  wire  m_567_io_in_1; // @[MUL.scala 124:19]
  wire  m_567_io_out_0; // @[MUL.scala 124:19]
  wire  m_567_io_out_1; // @[MUL.scala 124:19]
  wire  m_568_io_in_0; // @[MUL.scala 124:19]
  wire  m_568_io_in_1; // @[MUL.scala 124:19]
  wire  m_568_io_out_0; // @[MUL.scala 124:19]
  wire  m_568_io_out_1; // @[MUL.scala 124:19]
  wire  m_569_io_in_0; // @[MUL.scala 124:19]
  wire  m_569_io_in_1; // @[MUL.scala 124:19]
  wire  m_569_io_out_0; // @[MUL.scala 124:19]
  wire  m_569_io_out_1; // @[MUL.scala 124:19]
  wire  m_570_io_in_0; // @[MUL.scala 124:19]
  wire  m_570_io_in_1; // @[MUL.scala 124:19]
  wire  m_570_io_out_0; // @[MUL.scala 124:19]
  wire  m_570_io_out_1; // @[MUL.scala 124:19]
  wire  m_571_io_in_0; // @[MUL.scala 124:19]
  wire  m_571_io_in_1; // @[MUL.scala 124:19]
  wire  m_571_io_out_0; // @[MUL.scala 124:19]
  wire  m_571_io_out_1; // @[MUL.scala 124:19]
  wire  m_572_io_in_0; // @[MUL.scala 124:19]
  wire  m_572_io_in_1; // @[MUL.scala 124:19]
  wire  m_572_io_out_0; // @[MUL.scala 124:19]
  wire  m_572_io_out_1; // @[MUL.scala 124:19]
  wire  m_573_io_in_0; // @[MUL.scala 124:19]
  wire  m_573_io_in_1; // @[MUL.scala 124:19]
  wire  m_573_io_out_0; // @[MUL.scala 124:19]
  wire  m_573_io_out_1; // @[MUL.scala 124:19]
  wire  m_574_io_in_0; // @[MUL.scala 124:19]
  wire  m_574_io_in_1; // @[MUL.scala 124:19]
  wire  m_574_io_out_0; // @[MUL.scala 124:19]
  wire  m_574_io_out_1; // @[MUL.scala 124:19]
  wire  m_575_io_in_0; // @[MUL.scala 124:19]
  wire  m_575_io_in_1; // @[MUL.scala 124:19]
  wire  m_575_io_out_0; // @[MUL.scala 124:19]
  wire  m_575_io_out_1; // @[MUL.scala 124:19]
  wire  m_576_io_in_0; // @[MUL.scala 124:19]
  wire  m_576_io_in_1; // @[MUL.scala 124:19]
  wire  m_576_io_out_0; // @[MUL.scala 124:19]
  wire  m_576_io_out_1; // @[MUL.scala 124:19]
  wire  m_577_io_in_0; // @[MUL.scala 124:19]
  wire  m_577_io_in_1; // @[MUL.scala 124:19]
  wire  m_577_io_out_0; // @[MUL.scala 124:19]
  wire  m_577_io_out_1; // @[MUL.scala 124:19]
  wire  m_578_io_in_0; // @[MUL.scala 124:19]
  wire  m_578_io_in_1; // @[MUL.scala 124:19]
  wire  m_578_io_out_0; // @[MUL.scala 124:19]
  wire  m_578_io_out_1; // @[MUL.scala 124:19]
  wire  m_579_io_in_0; // @[MUL.scala 124:19]
  wire  m_579_io_in_1; // @[MUL.scala 124:19]
  wire  m_579_io_out_0; // @[MUL.scala 124:19]
  wire  m_579_io_out_1; // @[MUL.scala 124:19]
  wire  m_580_io_in_0; // @[MUL.scala 124:19]
  wire  m_580_io_in_1; // @[MUL.scala 124:19]
  wire  m_580_io_out_0; // @[MUL.scala 124:19]
  wire  m_580_io_out_1; // @[MUL.scala 124:19]
  wire  m_581_io_in_0; // @[MUL.scala 124:19]
  wire  m_581_io_in_1; // @[MUL.scala 124:19]
  wire  m_581_io_out_0; // @[MUL.scala 124:19]
  wire  m_581_io_out_1; // @[MUL.scala 124:19]
  wire  m_582_io_in_0; // @[MUL.scala 124:19]
  wire  m_582_io_in_1; // @[MUL.scala 124:19]
  wire  m_582_io_out_0; // @[MUL.scala 124:19]
  wire  m_582_io_out_1; // @[MUL.scala 124:19]
  wire  m_583_io_in_0; // @[MUL.scala 124:19]
  wire  m_583_io_in_1; // @[MUL.scala 124:19]
  wire  m_583_io_out_0; // @[MUL.scala 124:19]
  wire  m_583_io_out_1; // @[MUL.scala 124:19]
  wire  m_584_io_in_0; // @[MUL.scala 124:19]
  wire  m_584_io_in_1; // @[MUL.scala 124:19]
  wire  m_584_io_out_0; // @[MUL.scala 124:19]
  wire  m_584_io_out_1; // @[MUL.scala 124:19]
  wire  m_585_io_in_0; // @[MUL.scala 124:19]
  wire  m_585_io_in_1; // @[MUL.scala 124:19]
  wire  m_585_io_out_0; // @[MUL.scala 124:19]
  wire  m_585_io_out_1; // @[MUL.scala 124:19]
  wire  m_586_io_in_0; // @[MUL.scala 124:19]
  wire  m_586_io_in_1; // @[MUL.scala 124:19]
  wire  m_586_io_out_0; // @[MUL.scala 124:19]
  wire  m_586_io_out_1; // @[MUL.scala 124:19]
  wire  m_587_io_in_0; // @[MUL.scala 124:19]
  wire  m_587_io_in_1; // @[MUL.scala 124:19]
  wire  m_587_io_out_0; // @[MUL.scala 124:19]
  wire  m_587_io_out_1; // @[MUL.scala 124:19]
  wire  m_588_io_in_0; // @[MUL.scala 124:19]
  wire  m_588_io_in_1; // @[MUL.scala 124:19]
  wire  m_588_io_out_0; // @[MUL.scala 124:19]
  wire  m_588_io_out_1; // @[MUL.scala 124:19]
  wire  m_589_io_in_0; // @[MUL.scala 124:19]
  wire  m_589_io_in_1; // @[MUL.scala 124:19]
  wire  m_589_io_out_0; // @[MUL.scala 124:19]
  wire  m_589_io_out_1; // @[MUL.scala 124:19]
  wire  m_590_io_x1; // @[MUL.scala 102:19]
  wire  m_590_io_x2; // @[MUL.scala 102:19]
  wire  m_590_io_x3; // @[MUL.scala 102:19]
  wire  m_590_io_s; // @[MUL.scala 102:19]
  wire  m_590_io_cout; // @[MUL.scala 102:19]
  wire  m_591_io_x1; // @[MUL.scala 102:19]
  wire  m_591_io_x2; // @[MUL.scala 102:19]
  wire  m_591_io_x3; // @[MUL.scala 102:19]
  wire  m_591_io_s; // @[MUL.scala 102:19]
  wire  m_591_io_cout; // @[MUL.scala 102:19]
  wire  m_592_io_x1; // @[MUL.scala 102:19]
  wire  m_592_io_x2; // @[MUL.scala 102:19]
  wire  m_592_io_x3; // @[MUL.scala 102:19]
  wire  m_592_io_s; // @[MUL.scala 102:19]
  wire  m_592_io_cout; // @[MUL.scala 102:19]
  wire  m_593_io_x1; // @[MUL.scala 102:19]
  wire  m_593_io_x2; // @[MUL.scala 102:19]
  wire  m_593_io_x3; // @[MUL.scala 102:19]
  wire  m_593_io_s; // @[MUL.scala 102:19]
  wire  m_593_io_cout; // @[MUL.scala 102:19]
  wire  m_594_io_x1; // @[MUL.scala 102:19]
  wire  m_594_io_x2; // @[MUL.scala 102:19]
  wire  m_594_io_x3; // @[MUL.scala 102:19]
  wire  m_594_io_s; // @[MUL.scala 102:19]
  wire  m_594_io_cout; // @[MUL.scala 102:19]
  wire  m_595_io_x1; // @[MUL.scala 102:19]
  wire  m_595_io_x2; // @[MUL.scala 102:19]
  wire  m_595_io_x3; // @[MUL.scala 102:19]
  wire  m_595_io_s; // @[MUL.scala 102:19]
  wire  m_595_io_cout; // @[MUL.scala 102:19]
  wire  m_596_io_x1; // @[MUL.scala 102:19]
  wire  m_596_io_x2; // @[MUL.scala 102:19]
  wire  m_596_io_x3; // @[MUL.scala 102:19]
  wire  m_596_io_s; // @[MUL.scala 102:19]
  wire  m_596_io_cout; // @[MUL.scala 102:19]
  wire  m_597_io_x1; // @[MUL.scala 102:19]
  wire  m_597_io_x2; // @[MUL.scala 102:19]
  wire  m_597_io_x3; // @[MUL.scala 102:19]
  wire  m_597_io_s; // @[MUL.scala 102:19]
  wire  m_597_io_cout; // @[MUL.scala 102:19]
  wire  m_598_io_x1; // @[MUL.scala 102:19]
  wire  m_598_io_x2; // @[MUL.scala 102:19]
  wire  m_598_io_x3; // @[MUL.scala 102:19]
  wire  m_598_io_s; // @[MUL.scala 102:19]
  wire  m_598_io_cout; // @[MUL.scala 102:19]
  wire  m_599_io_x1; // @[MUL.scala 102:19]
  wire  m_599_io_x2; // @[MUL.scala 102:19]
  wire  m_599_io_x3; // @[MUL.scala 102:19]
  wire  m_599_io_s; // @[MUL.scala 102:19]
  wire  m_599_io_cout; // @[MUL.scala 102:19]
  wire  m_600_io_x1; // @[MUL.scala 102:19]
  wire  m_600_io_x2; // @[MUL.scala 102:19]
  wire  m_600_io_x3; // @[MUL.scala 102:19]
  wire  m_600_io_s; // @[MUL.scala 102:19]
  wire  m_600_io_cout; // @[MUL.scala 102:19]
  wire  m_601_io_x1; // @[MUL.scala 102:19]
  wire  m_601_io_x2; // @[MUL.scala 102:19]
  wire  m_601_io_x3; // @[MUL.scala 102:19]
  wire  m_601_io_s; // @[MUL.scala 102:19]
  wire  m_601_io_cout; // @[MUL.scala 102:19]
  wire  m_602_io_x1; // @[MUL.scala 102:19]
  wire  m_602_io_x2; // @[MUL.scala 102:19]
  wire  m_602_io_x3; // @[MUL.scala 102:19]
  wire  m_602_io_s; // @[MUL.scala 102:19]
  wire  m_602_io_cout; // @[MUL.scala 102:19]
  wire  m_603_io_x1; // @[MUL.scala 102:19]
  wire  m_603_io_x2; // @[MUL.scala 102:19]
  wire  m_603_io_x3; // @[MUL.scala 102:19]
  wire  m_603_io_s; // @[MUL.scala 102:19]
  wire  m_603_io_cout; // @[MUL.scala 102:19]
  wire  m_604_io_x1; // @[MUL.scala 102:19]
  wire  m_604_io_x2; // @[MUL.scala 102:19]
  wire  m_604_io_x3; // @[MUL.scala 102:19]
  wire  m_604_io_s; // @[MUL.scala 102:19]
  wire  m_604_io_cout; // @[MUL.scala 102:19]
  wire  m_605_io_x1; // @[MUL.scala 102:19]
  wire  m_605_io_x2; // @[MUL.scala 102:19]
  wire  m_605_io_x3; // @[MUL.scala 102:19]
  wire  m_605_io_s; // @[MUL.scala 102:19]
  wire  m_605_io_cout; // @[MUL.scala 102:19]
  wire  m_606_io_x1; // @[MUL.scala 102:19]
  wire  m_606_io_x2; // @[MUL.scala 102:19]
  wire  m_606_io_x3; // @[MUL.scala 102:19]
  wire  m_606_io_s; // @[MUL.scala 102:19]
  wire  m_606_io_cout; // @[MUL.scala 102:19]
  wire  m_607_io_x1; // @[MUL.scala 102:19]
  wire  m_607_io_x2; // @[MUL.scala 102:19]
  wire  m_607_io_x3; // @[MUL.scala 102:19]
  wire  m_607_io_s; // @[MUL.scala 102:19]
  wire  m_607_io_cout; // @[MUL.scala 102:19]
  wire  m_608_io_x1; // @[MUL.scala 102:19]
  wire  m_608_io_x2; // @[MUL.scala 102:19]
  wire  m_608_io_x3; // @[MUL.scala 102:19]
  wire  m_608_io_s; // @[MUL.scala 102:19]
  wire  m_608_io_cout; // @[MUL.scala 102:19]
  wire  m_609_io_x1; // @[MUL.scala 102:19]
  wire  m_609_io_x2; // @[MUL.scala 102:19]
  wire  m_609_io_x3; // @[MUL.scala 102:19]
  wire  m_609_io_s; // @[MUL.scala 102:19]
  wire  m_609_io_cout; // @[MUL.scala 102:19]
  wire  m_610_io_x1; // @[MUL.scala 102:19]
  wire  m_610_io_x2; // @[MUL.scala 102:19]
  wire  m_610_io_x3; // @[MUL.scala 102:19]
  wire  m_610_io_s; // @[MUL.scala 102:19]
  wire  m_610_io_cout; // @[MUL.scala 102:19]
  wire  m_611_io_x1; // @[MUL.scala 102:19]
  wire  m_611_io_x2; // @[MUL.scala 102:19]
  wire  m_611_io_x3; // @[MUL.scala 102:19]
  wire  m_611_io_s; // @[MUL.scala 102:19]
  wire  m_611_io_cout; // @[MUL.scala 102:19]
  wire  m_612_io_x1; // @[MUL.scala 102:19]
  wire  m_612_io_x2; // @[MUL.scala 102:19]
  wire  m_612_io_x3; // @[MUL.scala 102:19]
  wire  m_612_io_s; // @[MUL.scala 102:19]
  wire  m_612_io_cout; // @[MUL.scala 102:19]
  wire  m_613_io_x1; // @[MUL.scala 102:19]
  wire  m_613_io_x2; // @[MUL.scala 102:19]
  wire  m_613_io_x3; // @[MUL.scala 102:19]
  wire  m_613_io_s; // @[MUL.scala 102:19]
  wire  m_613_io_cout; // @[MUL.scala 102:19]
  wire  m_614_io_x1; // @[MUL.scala 102:19]
  wire  m_614_io_x2; // @[MUL.scala 102:19]
  wire  m_614_io_x3; // @[MUL.scala 102:19]
  wire  m_614_io_s; // @[MUL.scala 102:19]
  wire  m_614_io_cout; // @[MUL.scala 102:19]
  wire  m_615_io_x1; // @[MUL.scala 102:19]
  wire  m_615_io_x2; // @[MUL.scala 102:19]
  wire  m_615_io_x3; // @[MUL.scala 102:19]
  wire  m_615_io_s; // @[MUL.scala 102:19]
  wire  m_615_io_cout; // @[MUL.scala 102:19]
  wire  m_616_io_x1; // @[MUL.scala 102:19]
  wire  m_616_io_x2; // @[MUL.scala 102:19]
  wire  m_616_io_x3; // @[MUL.scala 102:19]
  wire  m_616_io_s; // @[MUL.scala 102:19]
  wire  m_616_io_cout; // @[MUL.scala 102:19]
  wire  m_617_io_x1; // @[MUL.scala 102:19]
  wire  m_617_io_x2; // @[MUL.scala 102:19]
  wire  m_617_io_x3; // @[MUL.scala 102:19]
  wire  m_617_io_s; // @[MUL.scala 102:19]
  wire  m_617_io_cout; // @[MUL.scala 102:19]
  wire  m_618_io_x1; // @[MUL.scala 102:19]
  wire  m_618_io_x2; // @[MUL.scala 102:19]
  wire  m_618_io_x3; // @[MUL.scala 102:19]
  wire  m_618_io_s; // @[MUL.scala 102:19]
  wire  m_618_io_cout; // @[MUL.scala 102:19]
  wire  m_619_io_x1; // @[MUL.scala 102:19]
  wire  m_619_io_x2; // @[MUL.scala 102:19]
  wire  m_619_io_x3; // @[MUL.scala 102:19]
  wire  m_619_io_s; // @[MUL.scala 102:19]
  wire  m_619_io_cout; // @[MUL.scala 102:19]
  wire  m_620_io_x1; // @[MUL.scala 102:19]
  wire  m_620_io_x2; // @[MUL.scala 102:19]
  wire  m_620_io_x3; // @[MUL.scala 102:19]
  wire  m_620_io_s; // @[MUL.scala 102:19]
  wire  m_620_io_cout; // @[MUL.scala 102:19]
  wire  m_621_io_x1; // @[MUL.scala 102:19]
  wire  m_621_io_x2; // @[MUL.scala 102:19]
  wire  m_621_io_x3; // @[MUL.scala 102:19]
  wire  m_621_io_s; // @[MUL.scala 102:19]
  wire  m_621_io_cout; // @[MUL.scala 102:19]
  wire  m_622_io_x1; // @[MUL.scala 102:19]
  wire  m_622_io_x2; // @[MUL.scala 102:19]
  wire  m_622_io_x3; // @[MUL.scala 102:19]
  wire  m_622_io_s; // @[MUL.scala 102:19]
  wire  m_622_io_cout; // @[MUL.scala 102:19]
  wire  m_623_io_x1; // @[MUL.scala 102:19]
  wire  m_623_io_x2; // @[MUL.scala 102:19]
  wire  m_623_io_x3; // @[MUL.scala 102:19]
  wire  m_623_io_s; // @[MUL.scala 102:19]
  wire  m_623_io_cout; // @[MUL.scala 102:19]
  wire  m_624_io_in_0; // @[MUL.scala 124:19]
  wire  m_624_io_in_1; // @[MUL.scala 124:19]
  wire  m_624_io_out_0; // @[MUL.scala 124:19]
  wire  m_624_io_out_1; // @[MUL.scala 124:19]
  wire  m_625_io_in_0; // @[MUL.scala 124:19]
  wire  m_625_io_in_1; // @[MUL.scala 124:19]
  wire  m_625_io_out_0; // @[MUL.scala 124:19]
  wire  m_625_io_out_1; // @[MUL.scala 124:19]
  wire  m_626_io_in_0; // @[MUL.scala 124:19]
  wire  m_626_io_in_1; // @[MUL.scala 124:19]
  wire  m_626_io_out_0; // @[MUL.scala 124:19]
  wire  m_626_io_out_1; // @[MUL.scala 124:19]
  wire  m_627_io_in_0; // @[MUL.scala 124:19]
  wire  m_627_io_in_1; // @[MUL.scala 124:19]
  wire  m_627_io_out_0; // @[MUL.scala 124:19]
  wire  m_627_io_out_1; // @[MUL.scala 124:19]
  wire  m_628_io_in_0; // @[MUL.scala 124:19]
  wire  m_628_io_in_1; // @[MUL.scala 124:19]
  wire  m_628_io_out_0; // @[MUL.scala 124:19]
  wire  m_628_io_out_1; // @[MUL.scala 124:19]
  wire  m_629_io_in_0; // @[MUL.scala 124:19]
  wire  m_629_io_in_1; // @[MUL.scala 124:19]
  wire  m_629_io_out_0; // @[MUL.scala 124:19]
  wire  m_629_io_out_1; // @[MUL.scala 124:19]
  wire  m_630_io_in_0; // @[MUL.scala 124:19]
  wire  m_630_io_in_1; // @[MUL.scala 124:19]
  wire  m_630_io_out_0; // @[MUL.scala 124:19]
  wire  m_630_io_out_1; // @[MUL.scala 124:19]
  wire  m_631_io_in_0; // @[MUL.scala 124:19]
  wire  m_631_io_in_1; // @[MUL.scala 124:19]
  wire  m_631_io_out_0; // @[MUL.scala 124:19]
  wire  m_631_io_out_1; // @[MUL.scala 124:19]
  wire  m_632_io_in_0; // @[MUL.scala 124:19]
  wire  m_632_io_in_1; // @[MUL.scala 124:19]
  wire  m_632_io_out_0; // @[MUL.scala 124:19]
  wire  m_632_io_out_1; // @[MUL.scala 124:19]
  wire  m_633_io_in_0; // @[MUL.scala 124:19]
  wire  m_633_io_in_1; // @[MUL.scala 124:19]
  wire  m_633_io_out_0; // @[MUL.scala 124:19]
  wire  m_633_io_out_1; // @[MUL.scala 124:19]
  wire  m_634_io_in_0; // @[MUL.scala 124:19]
  wire  m_634_io_in_1; // @[MUL.scala 124:19]
  wire  m_634_io_out_0; // @[MUL.scala 124:19]
  wire  m_634_io_out_1; // @[MUL.scala 124:19]
  wire  m_635_io_in_0; // @[MUL.scala 124:19]
  wire  m_635_io_in_1; // @[MUL.scala 124:19]
  wire  m_635_io_out_0; // @[MUL.scala 124:19]
  wire  m_635_io_out_1; // @[MUL.scala 124:19]
  wire  m_636_io_in_0; // @[MUL.scala 124:19]
  wire  m_636_io_in_1; // @[MUL.scala 124:19]
  wire  m_636_io_out_0; // @[MUL.scala 124:19]
  wire  m_636_io_out_1; // @[MUL.scala 124:19]
  wire  m_637_io_in_0; // @[MUL.scala 124:19]
  wire  m_637_io_in_1; // @[MUL.scala 124:19]
  wire  m_637_io_out_0; // @[MUL.scala 124:19]
  wire  m_637_io_out_1; // @[MUL.scala 124:19]
  wire  m_638_io_in_0; // @[MUL.scala 124:19]
  wire  m_638_io_in_1; // @[MUL.scala 124:19]
  wire  m_638_io_out_0; // @[MUL.scala 124:19]
  wire  m_638_io_out_1; // @[MUL.scala 124:19]
  wire  m_639_io_in_0; // @[MUL.scala 124:19]
  wire  m_639_io_in_1; // @[MUL.scala 124:19]
  wire  m_639_io_out_0; // @[MUL.scala 124:19]
  wire  m_639_io_out_1; // @[MUL.scala 124:19]
  wire  m_640_io_in_0; // @[MUL.scala 124:19]
  wire  m_640_io_in_1; // @[MUL.scala 124:19]
  wire  m_640_io_out_0; // @[MUL.scala 124:19]
  wire  m_640_io_out_1; // @[MUL.scala 124:19]
  wire  m_641_io_in_0; // @[MUL.scala 124:19]
  wire  m_641_io_in_1; // @[MUL.scala 124:19]
  wire  m_641_io_out_0; // @[MUL.scala 124:19]
  wire  m_641_io_out_1; // @[MUL.scala 124:19]
  wire  m_642_io_in_0; // @[MUL.scala 124:19]
  wire  m_642_io_in_1; // @[MUL.scala 124:19]
  wire  m_642_io_out_0; // @[MUL.scala 124:19]
  wire  m_642_io_out_1; // @[MUL.scala 124:19]
  wire  m_643_io_in_0; // @[MUL.scala 124:19]
  wire  m_643_io_in_1; // @[MUL.scala 124:19]
  wire  m_643_io_out_0; // @[MUL.scala 124:19]
  wire  m_643_io_out_1; // @[MUL.scala 124:19]
  wire  m_644_io_in_0; // @[MUL.scala 124:19]
  wire  m_644_io_in_1; // @[MUL.scala 124:19]
  wire  m_644_io_out_0; // @[MUL.scala 124:19]
  wire  m_644_io_out_1; // @[MUL.scala 124:19]
  wire  m_645_io_in_0; // @[MUL.scala 124:19]
  wire  m_645_io_in_1; // @[MUL.scala 124:19]
  wire  m_645_io_out_0; // @[MUL.scala 124:19]
  wire  m_645_io_out_1; // @[MUL.scala 124:19]
  wire  m_646_io_in_0; // @[MUL.scala 124:19]
  wire  m_646_io_in_1; // @[MUL.scala 124:19]
  wire  m_646_io_out_0; // @[MUL.scala 124:19]
  wire  m_646_io_out_1; // @[MUL.scala 124:19]
  wire  m_647_io_in_0; // @[MUL.scala 124:19]
  wire  m_647_io_in_1; // @[MUL.scala 124:19]
  wire  m_647_io_out_0; // @[MUL.scala 124:19]
  wire  m_647_io_out_1; // @[MUL.scala 124:19]
  wire  m_648_io_in_0; // @[MUL.scala 124:19]
  wire  m_648_io_in_1; // @[MUL.scala 124:19]
  wire  m_648_io_out_0; // @[MUL.scala 124:19]
  wire  m_648_io_out_1; // @[MUL.scala 124:19]
  wire  m_649_io_in_0; // @[MUL.scala 124:19]
  wire  m_649_io_in_1; // @[MUL.scala 124:19]
  wire  m_649_io_out_0; // @[MUL.scala 124:19]
  wire  m_649_io_out_1; // @[MUL.scala 124:19]
  wire  m_650_io_in_0; // @[MUL.scala 124:19]
  wire  m_650_io_in_1; // @[MUL.scala 124:19]
  wire  m_650_io_out_0; // @[MUL.scala 124:19]
  wire  m_650_io_out_1; // @[MUL.scala 124:19]
  wire  m_651_io_in_0; // @[MUL.scala 124:19]
  wire  m_651_io_in_1; // @[MUL.scala 124:19]
  wire  m_651_io_out_0; // @[MUL.scala 124:19]
  wire  m_651_io_out_1; // @[MUL.scala 124:19]
  wire  m_652_io_in_0; // @[MUL.scala 124:19]
  wire  m_652_io_in_1; // @[MUL.scala 124:19]
  wire  m_652_io_out_0; // @[MUL.scala 124:19]
  wire  m_652_io_out_1; // @[MUL.scala 124:19]
  wire  m_653_io_in_0; // @[MUL.scala 124:19]
  wire  m_653_io_in_1; // @[MUL.scala 124:19]
  wire  m_653_io_out_0; // @[MUL.scala 124:19]
  wire  m_653_io_out_1; // @[MUL.scala 124:19]
  wire  m_654_io_in_0; // @[MUL.scala 124:19]
  wire  m_654_io_in_1; // @[MUL.scala 124:19]
  wire  m_654_io_out_0; // @[MUL.scala 124:19]
  wire  m_654_io_out_1; // @[MUL.scala 124:19]
  wire  m_655_io_in_0; // @[MUL.scala 124:19]
  wire  m_655_io_in_1; // @[MUL.scala 124:19]
  wire  m_655_io_out_0; // @[MUL.scala 124:19]
  wire  m_655_io_out_1; // @[MUL.scala 124:19]
  wire  m_656_io_in_0; // @[MUL.scala 124:19]
  wire  m_656_io_in_1; // @[MUL.scala 124:19]
  wire  m_656_io_out_0; // @[MUL.scala 124:19]
  wire  m_656_io_out_1; // @[MUL.scala 124:19]
  wire  m_657_io_in_0; // @[MUL.scala 124:19]
  wire  m_657_io_in_1; // @[MUL.scala 124:19]
  wire  m_657_io_out_0; // @[MUL.scala 124:19]
  wire  m_657_io_out_1; // @[MUL.scala 124:19]
  wire  m_658_io_in_0; // @[MUL.scala 124:19]
  wire  m_658_io_in_1; // @[MUL.scala 124:19]
  wire  m_658_io_out_0; // @[MUL.scala 124:19]
  wire  m_658_io_out_1; // @[MUL.scala 124:19]
  wire  m_659_io_in_0; // @[MUL.scala 124:19]
  wire  m_659_io_in_1; // @[MUL.scala 124:19]
  wire  m_659_io_out_0; // @[MUL.scala 124:19]
  wire  m_659_io_out_1; // @[MUL.scala 124:19]
  wire  m_660_io_in_0; // @[MUL.scala 124:19]
  wire  m_660_io_in_1; // @[MUL.scala 124:19]
  wire  m_660_io_out_0; // @[MUL.scala 124:19]
  wire  m_660_io_out_1; // @[MUL.scala 124:19]
  wire  m_661_io_x1; // @[MUL.scala 102:19]
  wire  m_661_io_x2; // @[MUL.scala 102:19]
  wire  m_661_io_x3; // @[MUL.scala 102:19]
  wire  m_661_io_s; // @[MUL.scala 102:19]
  wire  m_661_io_cout; // @[MUL.scala 102:19]
  wire  m_662_io_x1; // @[MUL.scala 102:19]
  wire  m_662_io_x2; // @[MUL.scala 102:19]
  wire  m_662_io_x3; // @[MUL.scala 102:19]
  wire  m_662_io_s; // @[MUL.scala 102:19]
  wire  m_662_io_cout; // @[MUL.scala 102:19]
  wire  m_663_io_x1; // @[MUL.scala 102:19]
  wire  m_663_io_x2; // @[MUL.scala 102:19]
  wire  m_663_io_x3; // @[MUL.scala 102:19]
  wire  m_663_io_s; // @[MUL.scala 102:19]
  wire  m_663_io_cout; // @[MUL.scala 102:19]
  wire  m_664_io_x1; // @[MUL.scala 102:19]
  wire  m_664_io_x2; // @[MUL.scala 102:19]
  wire  m_664_io_x3; // @[MUL.scala 102:19]
  wire  m_664_io_s; // @[MUL.scala 102:19]
  wire  m_664_io_cout; // @[MUL.scala 102:19]
  wire  m_665_io_x1; // @[MUL.scala 102:19]
  wire  m_665_io_x2; // @[MUL.scala 102:19]
  wire  m_665_io_x3; // @[MUL.scala 102:19]
  wire  m_665_io_s; // @[MUL.scala 102:19]
  wire  m_665_io_cout; // @[MUL.scala 102:19]
  wire  m_666_io_x1; // @[MUL.scala 102:19]
  wire  m_666_io_x2; // @[MUL.scala 102:19]
  wire  m_666_io_x3; // @[MUL.scala 102:19]
  wire  m_666_io_s; // @[MUL.scala 102:19]
  wire  m_666_io_cout; // @[MUL.scala 102:19]
  wire  m_667_io_x1; // @[MUL.scala 102:19]
  wire  m_667_io_x2; // @[MUL.scala 102:19]
  wire  m_667_io_x3; // @[MUL.scala 102:19]
  wire  m_667_io_s; // @[MUL.scala 102:19]
  wire  m_667_io_cout; // @[MUL.scala 102:19]
  wire  m_668_io_x1; // @[MUL.scala 102:19]
  wire  m_668_io_x2; // @[MUL.scala 102:19]
  wire  m_668_io_x3; // @[MUL.scala 102:19]
  wire  m_668_io_s; // @[MUL.scala 102:19]
  wire  m_668_io_cout; // @[MUL.scala 102:19]
  wire  m_669_io_x1; // @[MUL.scala 102:19]
  wire  m_669_io_x2; // @[MUL.scala 102:19]
  wire  m_669_io_x3; // @[MUL.scala 102:19]
  wire  m_669_io_s; // @[MUL.scala 102:19]
  wire  m_669_io_cout; // @[MUL.scala 102:19]
  wire  m_670_io_x1; // @[MUL.scala 102:19]
  wire  m_670_io_x2; // @[MUL.scala 102:19]
  wire  m_670_io_x3; // @[MUL.scala 102:19]
  wire  m_670_io_s; // @[MUL.scala 102:19]
  wire  m_670_io_cout; // @[MUL.scala 102:19]
  wire  m_671_io_x1; // @[MUL.scala 102:19]
  wire  m_671_io_x2; // @[MUL.scala 102:19]
  wire  m_671_io_x3; // @[MUL.scala 102:19]
  wire  m_671_io_s; // @[MUL.scala 102:19]
  wire  m_671_io_cout; // @[MUL.scala 102:19]
  wire  m_672_io_x1; // @[MUL.scala 102:19]
  wire  m_672_io_x2; // @[MUL.scala 102:19]
  wire  m_672_io_x3; // @[MUL.scala 102:19]
  wire  m_672_io_s; // @[MUL.scala 102:19]
  wire  m_672_io_cout; // @[MUL.scala 102:19]
  wire  m_673_io_x1; // @[MUL.scala 102:19]
  wire  m_673_io_x2; // @[MUL.scala 102:19]
  wire  m_673_io_x3; // @[MUL.scala 102:19]
  wire  m_673_io_s; // @[MUL.scala 102:19]
  wire  m_673_io_cout; // @[MUL.scala 102:19]
  wire  m_674_io_x1; // @[MUL.scala 102:19]
  wire  m_674_io_x2; // @[MUL.scala 102:19]
  wire  m_674_io_x3; // @[MUL.scala 102:19]
  wire  m_674_io_s; // @[MUL.scala 102:19]
  wire  m_674_io_cout; // @[MUL.scala 102:19]
  wire  m_675_io_x1; // @[MUL.scala 102:19]
  wire  m_675_io_x2; // @[MUL.scala 102:19]
  wire  m_675_io_x3; // @[MUL.scala 102:19]
  wire  m_675_io_s; // @[MUL.scala 102:19]
  wire  m_675_io_cout; // @[MUL.scala 102:19]
  wire  m_676_io_x1; // @[MUL.scala 102:19]
  wire  m_676_io_x2; // @[MUL.scala 102:19]
  wire  m_676_io_x3; // @[MUL.scala 102:19]
  wire  m_676_io_s; // @[MUL.scala 102:19]
  wire  m_676_io_cout; // @[MUL.scala 102:19]
  wire  m_677_io_x1; // @[MUL.scala 102:19]
  wire  m_677_io_x2; // @[MUL.scala 102:19]
  wire  m_677_io_x3; // @[MUL.scala 102:19]
  wire  m_677_io_s; // @[MUL.scala 102:19]
  wire  m_677_io_cout; // @[MUL.scala 102:19]
  wire  m_678_io_x1; // @[MUL.scala 102:19]
  wire  m_678_io_x2; // @[MUL.scala 102:19]
  wire  m_678_io_x3; // @[MUL.scala 102:19]
  wire  m_678_io_s; // @[MUL.scala 102:19]
  wire  m_678_io_cout; // @[MUL.scala 102:19]
  wire  m_679_io_in_0; // @[MUL.scala 124:19]
  wire  m_679_io_in_1; // @[MUL.scala 124:19]
  wire  m_679_io_out_0; // @[MUL.scala 124:19]
  wire  m_679_io_out_1; // @[MUL.scala 124:19]
  wire  m_680_io_in_0; // @[MUL.scala 124:19]
  wire  m_680_io_in_1; // @[MUL.scala 124:19]
  wire  m_680_io_out_0; // @[MUL.scala 124:19]
  wire  m_680_io_out_1; // @[MUL.scala 124:19]
  wire  m_681_io_in_0; // @[MUL.scala 124:19]
  wire  m_681_io_in_1; // @[MUL.scala 124:19]
  wire  m_681_io_out_0; // @[MUL.scala 124:19]
  wire  m_681_io_out_1; // @[MUL.scala 124:19]
  wire  m_682_io_in_0; // @[MUL.scala 124:19]
  wire  m_682_io_in_1; // @[MUL.scala 124:19]
  wire  m_682_io_out_0; // @[MUL.scala 124:19]
  wire  m_682_io_out_1; // @[MUL.scala 124:19]
  wire  m_683_io_in_0; // @[MUL.scala 124:19]
  wire  m_683_io_in_1; // @[MUL.scala 124:19]
  wire  m_683_io_out_0; // @[MUL.scala 124:19]
  wire  m_683_io_out_1; // @[MUL.scala 124:19]
  wire  m_684_io_in_0; // @[MUL.scala 124:19]
  wire  m_684_io_in_1; // @[MUL.scala 124:19]
  wire  m_684_io_out_0; // @[MUL.scala 124:19]
  wire  m_684_io_out_1; // @[MUL.scala 124:19]
  wire  m_685_io_in_0; // @[MUL.scala 124:19]
  wire  m_685_io_in_1; // @[MUL.scala 124:19]
  wire  m_685_io_out_0; // @[MUL.scala 124:19]
  wire  m_685_io_out_1; // @[MUL.scala 124:19]
  wire  m_686_io_in_0; // @[MUL.scala 124:19]
  wire  m_686_io_in_1; // @[MUL.scala 124:19]
  wire  m_686_io_out_0; // @[MUL.scala 124:19]
  wire  m_686_io_out_1; // @[MUL.scala 124:19]
  wire  m_687_io_in_0; // @[MUL.scala 124:19]
  wire  m_687_io_in_1; // @[MUL.scala 124:19]
  wire  m_687_io_out_0; // @[MUL.scala 124:19]
  wire  m_687_io_out_1; // @[MUL.scala 124:19]
  wire  m_688_io_in_0; // @[MUL.scala 124:19]
  wire  m_688_io_in_1; // @[MUL.scala 124:19]
  wire  m_688_io_out_0; // @[MUL.scala 124:19]
  wire  m_688_io_out_1; // @[MUL.scala 124:19]
  wire  m_689_io_in_0; // @[MUL.scala 124:19]
  wire  m_689_io_in_1; // @[MUL.scala 124:19]
  wire  m_689_io_out_0; // @[MUL.scala 124:19]
  wire  m_689_io_out_1; // @[MUL.scala 124:19]
  wire  m_690_io_in_0; // @[MUL.scala 124:19]
  wire  m_690_io_in_1; // @[MUL.scala 124:19]
  wire  m_690_io_out_0; // @[MUL.scala 124:19]
  wire  m_690_io_out_1; // @[MUL.scala 124:19]
  wire  m_691_io_in_0; // @[MUL.scala 124:19]
  wire  m_691_io_in_1; // @[MUL.scala 124:19]
  wire  m_691_io_out_0; // @[MUL.scala 124:19]
  wire  m_691_io_out_1; // @[MUL.scala 124:19]
  wire  m_692_io_in_0; // @[MUL.scala 124:19]
  wire  m_692_io_in_1; // @[MUL.scala 124:19]
  wire  m_692_io_out_0; // @[MUL.scala 124:19]
  wire  m_692_io_out_1; // @[MUL.scala 124:19]
  wire  m_693_io_in_0; // @[MUL.scala 124:19]
  wire  m_693_io_in_1; // @[MUL.scala 124:19]
  wire  m_693_io_out_0; // @[MUL.scala 124:19]
  wire  m_693_io_out_1; // @[MUL.scala 124:19]
  wire  m_694_io_in_0; // @[MUL.scala 124:19]
  wire  m_694_io_in_1; // @[MUL.scala 124:19]
  wire  m_694_io_out_0; // @[MUL.scala 124:19]
  wire  m_694_io_out_1; // @[MUL.scala 124:19]
  wire  m_695_io_in_0; // @[MUL.scala 124:19]
  wire  m_695_io_in_1; // @[MUL.scala 124:19]
  wire  m_695_io_out_0; // @[MUL.scala 124:19]
  wire  m_695_io_out_1; // @[MUL.scala 124:19]
  wire  m_696_io_in_0; // @[MUL.scala 124:19]
  wire  m_696_io_in_1; // @[MUL.scala 124:19]
  wire  m_696_io_out_0; // @[MUL.scala 124:19]
  wire  m_696_io_out_1; // @[MUL.scala 124:19]
  wire  m_697_io_in_0; // @[MUL.scala 124:19]
  wire  m_697_io_in_1; // @[MUL.scala 124:19]
  wire  m_697_io_out_0; // @[MUL.scala 124:19]
  wire  m_697_io_out_1; // @[MUL.scala 124:19]
  wire  m_698_io_in_0; // @[MUL.scala 124:19]
  wire  m_698_io_in_1; // @[MUL.scala 124:19]
  wire  m_698_io_out_0; // @[MUL.scala 124:19]
  wire  m_698_io_out_1; // @[MUL.scala 124:19]
  wire  m_699_io_in_0; // @[MUL.scala 124:19]
  wire  m_699_io_in_1; // @[MUL.scala 124:19]
  wire  m_699_io_out_0; // @[MUL.scala 124:19]
  wire  m_699_io_out_1; // @[MUL.scala 124:19]
  wire  m_700_io_in_0; // @[MUL.scala 124:19]
  wire  m_700_io_in_1; // @[MUL.scala 124:19]
  wire  m_700_io_out_0; // @[MUL.scala 124:19]
  wire  m_700_io_out_1; // @[MUL.scala 124:19]
  wire  m_701_io_in_0; // @[MUL.scala 124:19]
  wire  m_701_io_in_1; // @[MUL.scala 124:19]
  wire  m_701_io_out_0; // @[MUL.scala 124:19]
  wire  m_701_io_out_1; // @[MUL.scala 124:19]
  wire  sign = io_in_bits_ctrl_data_src1[31]; // @[util.scala 11:19]
  wire [1:0] _T_1 = sign ? 2'h3 : 2'h0; // @[Bitwise.scala 77:12]
  wire [34:0] _T_3 = {_T_1,io_in_bits_ctrl_data_src1,1'h0}; // @[Cat.scala 33:92]
  wire  sign_1 = io_in_bits_ctrl_data_src2[31]; // @[util.scala 11:19]
  wire [1:0] _T_5 = sign_1 ? 2'h3 : 2'h0; // @[Bitwise.scala 77:12]
  wire [33:0] _T_6 = {_T_5,io_in_bits_ctrl_data_src2}; // @[Cat.scala 33:92]
  wire [33:0] _T_12 = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 33:92]
  wire [34:0] _T_15 = {2'h0,io_in_bits_ctrl_data_src1,1'h0}; // @[Cat.scala 33:92]
  wire  _src1_T = 2'h0 == io_in_bits_ctrl_flow_mul_sign; // @[util.scala 45:32]
  wire  _src1_T_1 = 2'h1 == io_in_bits_ctrl_flow_mul_sign; // @[util.scala 45:32]
  wire  _src1_T_2 = 2'h3 == io_in_bits_ctrl_flow_mul_sign; // @[util.scala 45:32]
  wire [34:0] _src1_T_3 = _src1_T ? _T_3 : 35'h0; // @[Mux.scala 27:73]
  wire [34:0] _src1_T_4 = _src1_T_1 ? _T_3 : 35'h0; // @[Mux.scala 27:73]
  wire [34:0] _src1_T_5 = _src1_T_2 ? _T_15 : 35'h0; // @[Mux.scala 27:73]
  wire [34:0] _src1_T_6 = _src1_T_3 | _src1_T_4; // @[Mux.scala 27:73]
  wire [34:0] src1 = _src1_T_6 | _src1_T_5; // @[Mux.scala 27:73]
  wire [33:0] _src2_T_3 = _src1_T ? _T_6 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _src2_T_4 = _src1_T_1 ? _T_12 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _src2_T_5 = _src1_T_2 ? _T_12 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _src2_T_6 = _src2_T_3 | _src2_T_4; // @[Mux.scala 27:73]
  wire  _T_56 = ~m_io_p[33]; // @[MUL.scala 323:93]
  wire  _T_93 = ~m_1_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_132 = ~m_2_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_171 = ~m_3_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_210 = ~m_4_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_249 = ~m_5_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_288 = ~m_6_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_327 = ~m_7_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_366 = ~m_8_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_405 = ~m_9_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_444 = ~m_10_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_483 = ~m_11_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_522 = ~m_12_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_561 = ~m_13_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_600 = ~m_14_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_639 = ~m_15_io_p[33]; // @[MUL.scala 317:92]
  wire  _T_678 = ~m_16_io_p[33]; // @[MUL.scala 326:92]
  reg  r; // @[Reg.scala 19:16]
  reg  r_1; // @[Reg.scala 19:16]
  reg  r_2; // @[Reg.scala 19:16]
  reg  r_3; // @[Reg.scala 19:16]
  reg  r_4; // @[Reg.scala 19:16]
  reg  r_5; // @[Reg.scala 19:16]
  reg  r_6; // @[Reg.scala 19:16]
  reg  r_7; // @[Reg.scala 19:16]
  reg  r_8; // @[Reg.scala 19:16]
  reg  r_9; // @[Reg.scala 19:16]
  reg  r_10; // @[Reg.scala 19:16]
  reg  r_11; // @[Reg.scala 19:16]
  reg  r_12; // @[Reg.scala 19:16]
  reg  r_13; // @[Reg.scala 19:16]
  reg  r_14; // @[Reg.scala 19:16]
  reg  r_15; // @[Reg.scala 19:16]
  reg  r_16; // @[Reg.scala 19:16]
  reg  r_17; // @[Reg.scala 19:16]
  reg  r_18; // @[Reg.scala 19:16]
  reg  r_19; // @[Reg.scala 19:16]
  reg  r_20; // @[Reg.scala 19:16]
  reg  r_21; // @[Reg.scala 19:16]
  reg  r_22; // @[Reg.scala 19:16]
  reg  r_23; // @[Reg.scala 19:16]
  reg  r_24; // @[Reg.scala 19:16]
  reg  r_25; // @[Reg.scala 19:16]
  reg  r_26; // @[Reg.scala 19:16]
  reg  r_27; // @[Reg.scala 19:16]
  reg  r_28; // @[Reg.scala 19:16]
  reg  r_29; // @[Reg.scala 19:16]
  reg  r_30; // @[Reg.scala 19:16]
  reg  r_31; // @[Reg.scala 19:16]
  reg  r_32; // @[Reg.scala 19:16]
  reg  r_33; // @[Reg.scala 19:16]
  reg  r_34; // @[Reg.scala 19:16]
  reg  r_35; // @[Reg.scala 19:16]
  reg  r_36; // @[Reg.scala 19:16]
  reg  r_37; // @[Reg.scala 19:16]
  reg  r_38; // @[Reg.scala 19:16]
  reg  r_39; // @[Reg.scala 19:16]
  reg  r_40; // @[Reg.scala 19:16]
  reg  r_41; // @[Reg.scala 19:16]
  reg  r_42; // @[Reg.scala 19:16]
  reg  r_43; // @[Reg.scala 19:16]
  reg  r_44; // @[Reg.scala 19:16]
  reg  r_45; // @[Reg.scala 19:16]
  reg  r_46; // @[Reg.scala 19:16]
  reg  r_47; // @[Reg.scala 19:16]
  reg  r_48; // @[Reg.scala 19:16]
  reg  r_49; // @[Reg.scala 19:16]
  reg  r_50; // @[Reg.scala 19:16]
  reg  r_51; // @[Reg.scala 19:16]
  reg  r_52; // @[Reg.scala 19:16]
  reg  r_53; // @[Reg.scala 19:16]
  reg  r_54; // @[Reg.scala 19:16]
  reg  r_55; // @[Reg.scala 19:16]
  reg  r_56; // @[Reg.scala 19:16]
  reg  r_57; // @[Reg.scala 19:16]
  reg  r_58; // @[Reg.scala 19:16]
  reg  r_59; // @[Reg.scala 19:16]
  reg  r_60; // @[Reg.scala 19:16]
  reg  r_61; // @[Reg.scala 19:16]
  reg  r_62; // @[Reg.scala 19:16]
  reg  r_63; // @[Reg.scala 19:16]
  reg  r_64; // @[Reg.scala 19:16]
  reg  r_65; // @[Reg.scala 19:16]
  reg  r_66; // @[Reg.scala 19:16]
  reg  r_67; // @[Reg.scala 19:16]
  reg  r_68; // @[Reg.scala 19:16]
  reg  r_69; // @[Reg.scala 19:16]
  reg  r_70; // @[Reg.scala 19:16]
  reg  r_71; // @[Reg.scala 19:16]
  reg  r_72; // @[Reg.scala 19:16]
  reg  r_73; // @[Reg.scala 19:16]
  reg  r_74; // @[Reg.scala 19:16]
  reg  r_75; // @[Reg.scala 19:16]
  reg  r_76; // @[Reg.scala 19:16]
  reg  r_77; // @[Reg.scala 19:16]
  reg  r_78; // @[Reg.scala 19:16]
  reg  r_79; // @[Reg.scala 19:16]
  reg  r_80; // @[Reg.scala 19:16]
  reg  r_81; // @[Reg.scala 19:16]
  reg  r_82; // @[Reg.scala 19:16]
  reg  r_83; // @[Reg.scala 19:16]
  reg  r_84; // @[Reg.scala 19:16]
  reg  r_85; // @[Reg.scala 19:16]
  reg  r_86; // @[Reg.scala 19:16]
  reg  r_87; // @[Reg.scala 19:16]
  reg  r_88; // @[Reg.scala 19:16]
  reg  r_89; // @[Reg.scala 19:16]
  reg  r_90; // @[Reg.scala 19:16]
  reg  r_91; // @[Reg.scala 19:16]
  reg  r_92; // @[Reg.scala 19:16]
  reg  r_93; // @[Reg.scala 19:16]
  reg  r_94; // @[Reg.scala 19:16]
  reg  r_95; // @[Reg.scala 19:16]
  reg  r_96; // @[Reg.scala 19:16]
  reg  r_97; // @[Reg.scala 19:16]
  reg  r_98; // @[Reg.scala 19:16]
  reg  r_99; // @[Reg.scala 19:16]
  reg  r_100; // @[Reg.scala 19:16]
  reg  r_101; // @[Reg.scala 19:16]
  reg  r_102; // @[Reg.scala 19:16]
  reg  r_103; // @[Reg.scala 19:16]
  reg  r_104; // @[Reg.scala 19:16]
  reg  r_105; // @[Reg.scala 19:16]
  reg  r_106; // @[Reg.scala 19:16]
  reg  r_107; // @[Reg.scala 19:16]
  reg  r_108; // @[Reg.scala 19:16]
  reg  r_109; // @[Reg.scala 19:16]
  reg  r_110; // @[Reg.scala 19:16]
  reg  r_111; // @[Reg.scala 19:16]
  reg  r_112; // @[Reg.scala 19:16]
  reg  r_113; // @[Reg.scala 19:16]
  reg  r_114; // @[Reg.scala 19:16]
  reg  r_115; // @[Reg.scala 19:16]
  reg  r_116; // @[Reg.scala 19:16]
  reg  r_117; // @[Reg.scala 19:16]
  reg  r_118; // @[Reg.scala 19:16]
  reg  r_119; // @[Reg.scala 19:16]
  reg  r_120; // @[Reg.scala 19:16]
  reg  r_121; // @[Reg.scala 19:16]
  reg  r_122; // @[Reg.scala 19:16]
  reg  r_123; // @[Reg.scala 19:16]
  reg  r_124; // @[Reg.scala 19:16]
  reg  r_125; // @[Reg.scala 19:16]
  reg  r_126; // @[Reg.scala 19:16]
  reg  r_127; // @[Reg.scala 19:16]
  reg  r_128; // @[Reg.scala 19:16]
  reg  r_129; // @[Reg.scala 19:16]
  reg  r_130; // @[Reg.scala 19:16]
  reg  r_131; // @[Reg.scala 19:16]
  reg  r_132; // @[Reg.scala 19:16]
  reg  r_133; // @[Reg.scala 19:16]
  reg  r_134; // @[Reg.scala 19:16]
  reg  r_135; // @[Reg.scala 19:16]
  reg  r_136; // @[Reg.scala 19:16]
  reg  r_137; // @[Reg.scala 19:16]
  reg  r_138; // @[Reg.scala 19:16]
  reg  r_139; // @[Reg.scala 19:16]
  reg  r_140; // @[Reg.scala 19:16]
  reg  r_141; // @[Reg.scala 19:16]
  reg  r_142; // @[Reg.scala 19:16]
  reg  r_143; // @[Reg.scala 19:16]
  reg  r_144; // @[Reg.scala 19:16]
  reg  r_145; // @[Reg.scala 19:16]
  reg  r_146; // @[Reg.scala 19:16]
  reg  r_147; // @[Reg.scala 19:16]
  reg  r_148; // @[Reg.scala 19:16]
  reg  r_149; // @[Reg.scala 19:16]
  reg  r_150; // @[Reg.scala 19:16]
  reg  r_151; // @[Reg.scala 19:16]
  reg  r_152; // @[Reg.scala 19:16]
  reg  r_153; // @[Reg.scala 19:16]
  reg  r_154; // @[Reg.scala 19:16]
  reg  r_155; // @[Reg.scala 19:16]
  reg  r_156; // @[Reg.scala 19:16]
  reg  r_157; // @[Reg.scala 19:16]
  reg  r_158; // @[Reg.scala 19:16]
  reg  r_159; // @[Reg.scala 19:16]
  reg  r_160; // @[Reg.scala 19:16]
  reg  r_161; // @[Reg.scala 19:16]
  reg  r_162; // @[Reg.scala 19:16]
  reg  r_163; // @[Reg.scala 19:16]
  reg  r_164; // @[Reg.scala 19:16]
  reg  r_165; // @[Reg.scala 19:16]
  reg  r_166; // @[Reg.scala 19:16]
  reg  r_167; // @[Reg.scala 19:16]
  reg  r_168; // @[Reg.scala 19:16]
  reg  r_169; // @[Reg.scala 19:16]
  reg  r_170; // @[Reg.scala 19:16]
  reg  r_171; // @[Reg.scala 19:16]
  reg  r_172; // @[Reg.scala 19:16]
  reg  r_173; // @[Reg.scala 19:16]
  reg  r_174; // @[Reg.scala 19:16]
  reg  r_175; // @[Reg.scala 19:16]
  reg  r_176; // @[Reg.scala 19:16]
  reg  r_177; // @[Reg.scala 19:16]
  reg  r_178; // @[Reg.scala 19:16]
  reg  r_179; // @[Reg.scala 19:16]
  reg  r_180; // @[Reg.scala 19:16]
  reg  r_181; // @[Reg.scala 19:16]
  reg  r_182; // @[Reg.scala 19:16]
  reg  r_183; // @[Reg.scala 19:16]
  reg  r_184; // @[Reg.scala 19:16]
  reg  r_185; // @[Reg.scala 19:16]
  reg  r_186; // @[Reg.scala 19:16]
  reg  r_187; // @[Reg.scala 19:16]
  reg  r_188; // @[Reg.scala 19:16]
  reg  r_189; // @[Reg.scala 19:16]
  reg  r_190; // @[Reg.scala 19:16]
  reg  r_191; // @[Reg.scala 19:16]
  reg  r_192; // @[Reg.scala 19:16]
  reg  r_193; // @[Reg.scala 19:16]
  reg  r_194; // @[Reg.scala 19:16]
  reg  r_195; // @[Reg.scala 19:16]
  reg  r_196; // @[Reg.scala 19:16]
  reg  r_197; // @[Reg.scala 19:16]
  reg  r_198; // @[Reg.scala 19:16]
  reg  r_199; // @[Reg.scala 19:16]
  reg  r_200; // @[Reg.scala 19:16]
  reg  r_201; // @[Reg.scala 19:16]
  reg  r_202; // @[Reg.scala 19:16]
  reg  r_203; // @[Reg.scala 19:16]
  reg  r_204; // @[Reg.scala 19:16]
  reg  r_205; // @[Reg.scala 19:16]
  reg  r_206; // @[Reg.scala 19:16]
  reg  r_207; // @[Reg.scala 19:16]
  reg  r_208; // @[Reg.scala 19:16]
  reg  r_209; // @[Reg.scala 19:16]
  reg  r_210; // @[Reg.scala 19:16]
  reg  r_211; // @[Reg.scala 19:16]
  reg  r_212; // @[Reg.scala 19:16]
  reg  r_213; // @[Reg.scala 19:16]
  reg  r_214; // @[Reg.scala 19:16]
  reg  r_215; // @[Reg.scala 19:16]
  reg  r_216; // @[Reg.scala 19:16]
  reg  r_217; // @[Reg.scala 19:16]
  reg  r_218; // @[Reg.scala 19:16]
  reg  r_219; // @[Reg.scala 19:16]
  reg  r_220; // @[Reg.scala 19:16]
  reg  r_221; // @[Reg.scala 19:16]
  reg  r_222; // @[Reg.scala 19:16]
  reg  r_223; // @[Reg.scala 19:16]
  reg  r_224; // @[Reg.scala 19:16]
  reg  r_225; // @[Reg.scala 19:16]
  reg  r_226; // @[Reg.scala 19:16]
  reg  r_227; // @[Reg.scala 19:16]
  reg  r_228; // @[Reg.scala 19:16]
  reg  r_229; // @[Reg.scala 19:16]
  reg  r_230; // @[Reg.scala 19:16]
  reg  r_231; // @[Reg.scala 19:16]
  reg  r_232; // @[Reg.scala 19:16]
  reg  r_233; // @[Reg.scala 19:16]
  reg  r_234; // @[Reg.scala 19:16]
  reg  r_235; // @[Reg.scala 19:16]
  reg  r_236; // @[Reg.scala 19:16]
  reg  r_237; // @[Reg.scala 19:16]
  reg  r_238; // @[Reg.scala 19:16]
  reg  r_239; // @[Reg.scala 19:16]
  reg  r_240; // @[Reg.scala 19:16]
  reg  r_241; // @[Reg.scala 19:16]
  reg  r_242; // @[Reg.scala 19:16]
  reg  r_243; // @[Reg.scala 19:16]
  reg  r_244; // @[Reg.scala 19:16]
  reg  r_245; // @[Reg.scala 19:16]
  reg  r_246; // @[Reg.scala 19:16]
  reg  r_247; // @[Reg.scala 19:16]
  reg  r_248; // @[Reg.scala 19:16]
  reg  r_249; // @[Reg.scala 19:16]
  reg  r_250; // @[Reg.scala 19:16]
  reg  r_251; // @[Reg.scala 19:16]
  reg  r_252; // @[Reg.scala 19:16]
  reg  r_253; // @[Reg.scala 19:16]
  reg  r_254; // @[Reg.scala 19:16]
  reg  r_255; // @[Reg.scala 19:16]
  reg  r_256; // @[Reg.scala 19:16]
  reg  r_257; // @[Reg.scala 19:16]
  reg  r_258; // @[Reg.scala 19:16]
  reg  r_259; // @[Reg.scala 19:16]
  reg  r_260; // @[Reg.scala 19:16]
  reg  r_261; // @[Reg.scala 19:16]
  reg  r_262; // @[Reg.scala 19:16]
  reg  r_263; // @[Reg.scala 19:16]
  reg  r_264; // @[Reg.scala 19:16]
  reg  r_265; // @[Reg.scala 19:16]
  reg  r_266; // @[Reg.scala 19:16]
  reg  r_267; // @[Reg.scala 19:16]
  reg  r_268; // @[Reg.scala 19:16]
  reg  r_269; // @[Reg.scala 19:16]
  reg  r_270; // @[Reg.scala 19:16]
  reg  r_271; // @[Reg.scala 19:16]
  reg  r_272; // @[Reg.scala 19:16]
  reg  r_273; // @[Reg.scala 19:16]
  reg  r_274; // @[Reg.scala 19:16]
  reg  r_275; // @[Reg.scala 19:16]
  reg  r_276; // @[Reg.scala 19:16]
  reg  r_277; // @[Reg.scala 19:16]
  reg  r_278; // @[Reg.scala 19:16]
  reg  r_279; // @[Reg.scala 19:16]
  reg  r_280; // @[Reg.scala 19:16]
  reg  r_281; // @[Reg.scala 19:16]
  reg  r_282; // @[Reg.scala 19:16]
  reg  r_283; // @[Reg.scala 19:16]
  reg  r_284; // @[Reg.scala 19:16]
  reg  r_285; // @[Reg.scala 19:16]
  reg  r_286; // @[Reg.scala 19:16]
  reg  r_287; // @[Reg.scala 19:16]
  reg  r_288; // @[Reg.scala 19:16]
  reg  r_289; // @[Reg.scala 19:16]
  reg  r_290; // @[Reg.scala 19:16]
  reg  r_291; // @[Reg.scala 19:16]
  reg  r_292; // @[Reg.scala 19:16]
  reg  r_293; // @[Reg.scala 19:16]
  reg  r_294; // @[Reg.scala 19:16]
  reg  r_295; // @[Reg.scala 19:16]
  reg  r_296; // @[Reg.scala 19:16]
  reg  r_297; // @[Reg.scala 19:16]
  reg  r_298; // @[Reg.scala 19:16]
  reg  r_299; // @[Reg.scala 19:16]
  reg  r_300; // @[Reg.scala 19:16]
  reg  r_301; // @[Reg.scala 19:16]
  reg  r_302; // @[Reg.scala 19:16]
  reg  r_303; // @[Reg.scala 19:16]
  reg  r_304; // @[Reg.scala 19:16]
  reg  r_305; // @[Reg.scala 19:16]
  reg  r_306; // @[Reg.scala 19:16]
  reg  r_307; // @[Reg.scala 19:16]
  reg  r_308; // @[Reg.scala 19:16]
  reg  r_309; // @[Reg.scala 19:16]
  reg  r_310; // @[Reg.scala 19:16]
  reg  r_311; // @[Reg.scala 19:16]
  reg  r_312; // @[Reg.scala 19:16]
  reg  r_313; // @[Reg.scala 19:16]
  reg  r_314; // @[Reg.scala 19:16]
  reg  r_315; // @[Reg.scala 19:16]
  reg  r_316; // @[Reg.scala 19:16]
  reg  r_317; // @[Reg.scala 19:16]
  reg  r_318; // @[Reg.scala 19:16]
  reg  r_319; // @[Reg.scala 19:16]
  reg  r_320; // @[Reg.scala 19:16]
  reg  r_321; // @[Reg.scala 19:16]
  reg  r_322; // @[Reg.scala 19:16]
  reg  r_323; // @[Reg.scala 19:16]
  reg  r_324; // @[Reg.scala 19:16]
  reg  r_325; // @[Reg.scala 19:16]
  reg  r_326; // @[Reg.scala 19:16]
  reg  r_327; // @[Reg.scala 19:16]
  reg  r_328; // @[Reg.scala 19:16]
  reg  r_329; // @[Reg.scala 19:16]
  reg  r_330; // @[Reg.scala 19:16]
  reg  r_331; // @[Reg.scala 19:16]
  reg  r_332; // @[Reg.scala 19:16]
  reg  r_333; // @[Reg.scala 19:16]
  reg  r_334; // @[Reg.scala 19:16]
  reg  r_335; // @[Reg.scala 19:16]
  reg  r_336; // @[Reg.scala 19:16]
  reg  r_337; // @[Reg.scala 19:16]
  reg  r_338; // @[Reg.scala 19:16]
  reg  r_339; // @[Reg.scala 19:16]
  reg  r_340; // @[Reg.scala 19:16]
  reg  r_341; // @[Reg.scala 19:16]
  reg  r_342; // @[Reg.scala 19:16]
  reg  r_343; // @[Reg.scala 19:16]
  reg  r_344; // @[Reg.scala 19:16]
  reg  r_345; // @[Reg.scala 19:16]
  reg  r_346; // @[Reg.scala 19:16]
  reg  r_347; // @[Reg.scala 19:16]
  reg  r_348; // @[Reg.scala 19:16]
  reg  r_349; // @[Reg.scala 19:16]
  reg  r_350; // @[Reg.scala 19:16]
  reg  r_351; // @[Reg.scala 19:16]
  reg  r_352; // @[Reg.scala 19:16]
  reg  r_353; // @[Reg.scala 19:16]
  reg  r_354; // @[Reg.scala 19:16]
  reg  r_355; // @[Reg.scala 19:16]
  reg  r_356; // @[Reg.scala 19:16]
  reg  r_357; // @[Reg.scala 19:16]
  reg  r_358; // @[Reg.scala 19:16]
  reg  r_359; // @[Reg.scala 19:16]
  reg  r_360; // @[Reg.scala 19:16]
  reg  r_361; // @[Reg.scala 19:16]
  reg  r_362; // @[Reg.scala 19:16]
  reg  r_363; // @[Reg.scala 19:16]
  reg  r_364; // @[Reg.scala 19:16]
  reg  r_365; // @[Reg.scala 19:16]
  reg  r_366; // @[Reg.scala 19:16]
  reg  r_367; // @[Reg.scala 19:16]
  reg  r_368; // @[Reg.scala 19:16]
  reg  r_369; // @[Reg.scala 19:16]
  reg  r_370; // @[Reg.scala 19:16]
  reg  r_371; // @[Reg.scala 19:16]
  reg  r_372; // @[Reg.scala 19:16]
  reg  r_373; // @[Reg.scala 19:16]
  reg  r_374; // @[Reg.scala 19:16]
  reg  r_375; // @[Reg.scala 19:16]
  reg  r_376; // @[Reg.scala 19:16]
  reg  r_377; // @[Reg.scala 19:16]
  reg  r_378; // @[Reg.scala 19:16]
  reg  r_379; // @[Reg.scala 19:16]
  reg  r_380; // @[Reg.scala 19:16]
  reg  r_381; // @[Reg.scala 19:16]
  reg  r_382; // @[Reg.scala 19:16]
  reg  r_383; // @[Reg.scala 19:16]
  reg  r_384; // @[Reg.scala 19:16]
  reg  r_385; // @[Reg.scala 19:16]
  reg  r_386; // @[Reg.scala 19:16]
  reg  r_387; // @[Reg.scala 19:16]
  reg  r_388; // @[Reg.scala 19:16]
  reg  r_390; // @[Reg.scala 19:16]
  reg  r_391; // @[Reg.scala 19:16]
  reg  r_392; // @[Reg.scala 19:16]
  reg  r_393; // @[Reg.scala 19:16]
  reg  r_394; // @[Reg.scala 19:16]
  reg  r_395; // @[Reg.scala 19:16]
  reg  r_396; // @[Reg.scala 19:16]
  reg  r_397; // @[Reg.scala 19:16]
  reg  r_398; // @[Reg.scala 19:16]
  reg  r_399; // @[Reg.scala 19:16]
  reg  r_400; // @[Reg.scala 19:16]
  reg  r_401; // @[Reg.scala 19:16]
  reg  r_402; // @[Reg.scala 19:16]
  reg  r_403; // @[Reg.scala 19:16]
  reg  r_404; // @[Reg.scala 19:16]
  reg  r_405; // @[Reg.scala 19:16]
  reg  r_406; // @[Reg.scala 19:16]
  reg  r_407; // @[Reg.scala 19:16]
  reg  r_408; // @[Reg.scala 19:16]
  reg  r_409; // @[Reg.scala 19:16]
  reg  r_410; // @[Reg.scala 19:16]
  reg  r_411; // @[Reg.scala 19:16]
  reg  r_412; // @[Reg.scala 19:16]
  reg  r_413; // @[Reg.scala 19:16]
  reg  r_414; // @[Reg.scala 19:16]
  reg  r_415; // @[Reg.scala 19:16]
  reg  r_416; // @[Reg.scala 19:16]
  reg  r_417; // @[Reg.scala 19:16]
  reg  r_418; // @[Reg.scala 19:16]
  reg  r_419; // @[Reg.scala 19:16]
  reg  r_421; // @[Reg.scala 19:16]
  reg  r_422; // @[Reg.scala 19:16]
  reg  r_423; // @[Reg.scala 19:16]
  reg  r_424; // @[Reg.scala 19:16]
  reg  r_425; // @[Reg.scala 19:16]
  reg  r_426; // @[Reg.scala 19:16]
  reg  r_427; // @[Reg.scala 19:16]
  reg  r_428; // @[Reg.scala 19:16]
  reg  r_429; // @[Reg.scala 19:16]
  reg  r_430; // @[Reg.scala 19:16]
  reg  r_431; // @[Reg.scala 19:16]
  reg  r_432; // @[Reg.scala 19:16]
  reg  r_433; // @[Reg.scala 19:16]
  reg  r_434; // @[Reg.scala 19:16]
  reg  r_435; // @[Reg.scala 19:16]
  reg  r_436; // @[Reg.scala 19:16]
  reg  r_437; // @[Reg.scala 19:16]
  reg  r_438; // @[Reg.scala 19:16]
  reg  r_439; // @[Reg.scala 19:16]
  reg  r_440; // @[Reg.scala 19:16]
  reg  r_441; // @[Reg.scala 19:16]
  reg  r_442; // @[Reg.scala 19:16]
  reg  r_443; // @[Reg.scala 19:16]
  reg  r_444; // @[Reg.scala 19:16]
  reg  r_445; // @[Reg.scala 19:16]
  reg  r_446; // @[Reg.scala 19:16]
  reg  r_447; // @[Reg.scala 19:16]
  reg  r_448; // @[Reg.scala 19:16]
  reg  r_450; // @[Reg.scala 19:16]
  reg  r_451; // @[Reg.scala 19:16]
  reg  r_452; // @[Reg.scala 19:16]
  reg  r_453; // @[Reg.scala 19:16]
  reg  r_454; // @[Reg.scala 19:16]
  reg  r_455; // @[Reg.scala 19:16]
  reg  r_456; // @[Reg.scala 19:16]
  reg  r_457; // @[Reg.scala 19:16]
  reg  r_458; // @[Reg.scala 19:16]
  reg  r_459; // @[Reg.scala 19:16]
  reg  r_460; // @[Reg.scala 19:16]
  reg  r_461; // @[Reg.scala 19:16]
  reg  r_462; // @[Reg.scala 19:16]
  reg  r_463; // @[Reg.scala 19:16]
  reg  r_464; // @[Reg.scala 19:16]
  reg  r_465; // @[Reg.scala 19:16]
  reg  r_466; // @[Reg.scala 19:16]
  reg  r_467; // @[Reg.scala 19:16]
  reg  r_468; // @[Reg.scala 19:16]
  reg  r_469; // @[Reg.scala 19:16]
  reg  r_470; // @[Reg.scala 19:16]
  reg  r_471; // @[Reg.scala 19:16]
  reg  r_472; // @[Reg.scala 19:16]
  reg  r_473; // @[Reg.scala 19:16]
  reg  r_474; // @[Reg.scala 19:16]
  reg  r_475; // @[Reg.scala 19:16]
  reg  r_477; // @[Reg.scala 19:16]
  reg  r_478; // @[Reg.scala 19:16]
  reg  r_479; // @[Reg.scala 19:16]
  reg  r_480; // @[Reg.scala 19:16]
  reg  r_481; // @[Reg.scala 19:16]
  reg  r_482; // @[Reg.scala 19:16]
  reg  r_483; // @[Reg.scala 19:16]
  reg  r_484; // @[Reg.scala 19:16]
  reg  r_485; // @[Reg.scala 19:16]
  reg  r_486; // @[Reg.scala 19:16]
  reg  r_487; // @[Reg.scala 19:16]
  reg  r_488; // @[Reg.scala 19:16]
  reg  r_489; // @[Reg.scala 19:16]
  reg  r_490; // @[Reg.scala 19:16]
  reg  r_491; // @[Reg.scala 19:16]
  reg  r_492; // @[Reg.scala 19:16]
  reg  r_493; // @[Reg.scala 19:16]
  reg  r_494; // @[Reg.scala 19:16]
  reg  r_495; // @[Reg.scala 19:16]
  reg  r_496; // @[Reg.scala 19:16]
  reg  r_497; // @[Reg.scala 19:16]
  reg  r_498; // @[Reg.scala 19:16]
  reg  r_499; // @[Reg.scala 19:16]
  reg  r_500; // @[Reg.scala 19:16]
  reg  r_502; // @[Reg.scala 19:16]
  reg  r_503; // @[Reg.scala 19:16]
  reg  r_504; // @[Reg.scala 19:16]
  reg  r_505; // @[Reg.scala 19:16]
  reg  r_506; // @[Reg.scala 19:16]
  reg  r_507; // @[Reg.scala 19:16]
  reg  r_508; // @[Reg.scala 19:16]
  reg  r_509; // @[Reg.scala 19:16]
  reg  r_510; // @[Reg.scala 19:16]
  reg  r_511; // @[Reg.scala 19:16]
  reg  r_512; // @[Reg.scala 19:16]
  reg  r_513; // @[Reg.scala 19:16]
  reg  r_514; // @[Reg.scala 19:16]
  reg  r_515; // @[Reg.scala 19:16]
  reg  r_516; // @[Reg.scala 19:16]
  reg  r_517; // @[Reg.scala 19:16]
  reg  r_518; // @[Reg.scala 19:16]
  reg  r_519; // @[Reg.scala 19:16]
  reg  r_520; // @[Reg.scala 19:16]
  reg  r_521; // @[Reg.scala 19:16]
  reg  r_522; // @[Reg.scala 19:16]
  reg  r_523; // @[Reg.scala 19:16]
  reg  r_525; // @[Reg.scala 19:16]
  reg  r_526; // @[Reg.scala 19:16]
  reg  r_527; // @[Reg.scala 19:16]
  reg  r_528; // @[Reg.scala 19:16]
  reg  r_529; // @[Reg.scala 19:16]
  reg  r_530; // @[Reg.scala 19:16]
  reg  r_531; // @[Reg.scala 19:16]
  reg  r_532; // @[Reg.scala 19:16]
  reg  r_533; // @[Reg.scala 19:16]
  reg  r_534; // @[Reg.scala 19:16]
  reg  r_535; // @[Reg.scala 19:16]
  reg  r_536; // @[Reg.scala 19:16]
  reg  r_537; // @[Reg.scala 19:16]
  reg  r_538; // @[Reg.scala 19:16]
  reg  r_539; // @[Reg.scala 19:16]
  reg  r_540; // @[Reg.scala 19:16]
  reg  r_541; // @[Reg.scala 19:16]
  reg  r_542; // @[Reg.scala 19:16]
  reg  r_543; // @[Reg.scala 19:16]
  reg  r_544; // @[Reg.scala 19:16]
  reg  r_546; // @[Reg.scala 19:16]
  reg  r_547; // @[Reg.scala 19:16]
  reg  r_548; // @[Reg.scala 19:16]
  reg  r_549; // @[Reg.scala 19:16]
  reg  r_550; // @[Reg.scala 19:16]
  reg  r_551; // @[Reg.scala 19:16]
  reg  r_552; // @[Reg.scala 19:16]
  reg  r_553; // @[Reg.scala 19:16]
  reg  r_554; // @[Reg.scala 19:16]
  reg  r_555; // @[Reg.scala 19:16]
  reg  r_556; // @[Reg.scala 19:16]
  reg  r_557; // @[Reg.scala 19:16]
  reg  r_558; // @[Reg.scala 19:16]
  reg  r_559; // @[Reg.scala 19:16]
  reg  r_560; // @[Reg.scala 19:16]
  reg  r_561; // @[Reg.scala 19:16]
  reg  r_562; // @[Reg.scala 19:16]
  reg  r_563; // @[Reg.scala 19:16]
  reg  r_565; // @[Reg.scala 19:16]
  reg  r_566; // @[Reg.scala 19:16]
  reg  r_567; // @[Reg.scala 19:16]
  reg  r_568; // @[Reg.scala 19:16]
  reg  r_569; // @[Reg.scala 19:16]
  reg  r_570; // @[Reg.scala 19:16]
  reg  r_571; // @[Reg.scala 19:16]
  reg  r_572; // @[Reg.scala 19:16]
  reg  r_573; // @[Reg.scala 19:16]
  reg  r_574; // @[Reg.scala 19:16]
  reg  r_575; // @[Reg.scala 19:16]
  reg  r_576; // @[Reg.scala 19:16]
  reg  r_577; // @[Reg.scala 19:16]
  reg  r_578; // @[Reg.scala 19:16]
  reg  r_579; // @[Reg.scala 19:16]
  reg  r_580; // @[Reg.scala 19:16]
  reg  r_582; // @[Reg.scala 19:16]
  reg  r_583; // @[Reg.scala 19:16]
  reg  r_584; // @[Reg.scala 19:16]
  reg  r_585; // @[Reg.scala 19:16]
  reg  r_586; // @[Reg.scala 19:16]
  reg  r_587; // @[Reg.scala 19:16]
  reg  r_588; // @[Reg.scala 19:16]
  reg  r_589; // @[Reg.scala 19:16]
  reg  r_590; // @[Reg.scala 19:16]
  reg  r_591; // @[Reg.scala 19:16]
  reg  r_592; // @[Reg.scala 19:16]
  reg  r_593; // @[Reg.scala 19:16]
  reg  r_594; // @[Reg.scala 19:16]
  reg  r_595; // @[Reg.scala 19:16]
  reg  r_597; // @[Reg.scala 19:16]
  reg  r_598; // @[Reg.scala 19:16]
  reg  r_599; // @[Reg.scala 19:16]
  reg  r_600; // @[Reg.scala 19:16]
  reg  r_601; // @[Reg.scala 19:16]
  reg  r_602; // @[Reg.scala 19:16]
  reg  r_603; // @[Reg.scala 19:16]
  reg  r_604; // @[Reg.scala 19:16]
  reg  r_605; // @[Reg.scala 19:16]
  reg  r_606; // @[Reg.scala 19:16]
  reg  r_607; // @[Reg.scala 19:16]
  reg  r_608; // @[Reg.scala 19:16]
  reg  r_610; // @[Reg.scala 19:16]
  reg  r_611; // @[Reg.scala 19:16]
  reg  r_612; // @[Reg.scala 19:16]
  reg  r_613; // @[Reg.scala 19:16]
  reg  r_614; // @[Reg.scala 19:16]
  reg  r_615; // @[Reg.scala 19:16]
  reg  r_616; // @[Reg.scala 19:16]
  reg  r_617; // @[Reg.scala 19:16]
  reg  r_618; // @[Reg.scala 19:16]
  reg  r_619; // @[Reg.scala 19:16]
  reg  r_621; // @[Reg.scala 19:16]
  reg  r_622; // @[Reg.scala 19:16]
  reg  r_623; // @[Reg.scala 19:16]
  reg  r_624; // @[Reg.scala 19:16]
  reg  r_625; // @[Reg.scala 19:16]
  reg  r_626; // @[Reg.scala 19:16]
  reg  r_627; // @[Reg.scala 19:16]
  reg  r_628; // @[Reg.scala 19:16]
  reg  r_630; // @[Reg.scala 19:16]
  reg  r_631; // @[Reg.scala 19:16]
  reg  r_632; // @[Reg.scala 19:16]
  reg  r_633; // @[Reg.scala 19:16]
  reg  r_634; // @[Reg.scala 19:16]
  reg  r_635; // @[Reg.scala 19:16]
  reg  r_637; // @[Reg.scala 19:16]
  reg  r_638; // @[Reg.scala 19:16]
  reg  r_639; // @[Reg.scala 19:16]
  reg  r_640; // @[Reg.scala 19:16]
  reg  r_642; // @[Reg.scala 19:16]
  reg  r_643; // @[Reg.scala 19:16]
  wire  c_1_92 = m_409_io_cout; // @[MUL.scala 263:22]
  wire  c_1_93 = m_411_io_cout; // @[MUL.scala 263:22]
  wire  c_1_94 = m_413_io_cout; // @[MUL.scala 263:22]
  wire  c_1_95 = m_415_io_cout; // @[MUL.scala 263:22]
  wire  c_1_114 = m_463_io_cout; // @[MUL.scala 263:22]
  wire  c_1_115 = m_465_io_cout; // @[MUL.scala 263:22]
  wire  c_1_116 = m_467_io_cout; // @[MUL.scala 263:22]
  wire  c_1_117 = m_469_io_cout; // @[MUL.scala 263:22]
  wire  c_1_118 = m_471_io_cout; // @[MUL.scala 263:22]
  wire  c_1_119 = m_473_io_cout; // @[MUL.scala 263:22]
  wire  c_1_120 = m_475_io_cout; // @[MUL.scala 263:22]
  wire  c_1_121 = m_477_io_cout; // @[MUL.scala 263:22]
  wire  s_0_174 = m_503_io_s; // @[MUL.scala 262:21]
  wire  c_0_174 = m_503_io_cout; // @[MUL.scala 263:22]
  wire  s_0_175 = m_504_io_s; // @[MUL.scala 262:21]
  wire  c_0_175 = m_504_io_cout; // @[MUL.scala 263:22]
  wire  s_0_176 = m_505_io_s; // @[MUL.scala 262:21]
  wire  c_0_176 = m_505_io_cout; // @[MUL.scala 263:22]
  wire  s_0_177 = m_506_io_s; // @[MUL.scala 262:21]
  wire  c_0_177 = m_506_io_cout; // @[MUL.scala 263:22]
  wire  s_0_178 = m_507_io_s; // @[MUL.scala 262:21]
  wire  c_0_178 = m_507_io_cout; // @[MUL.scala 263:22]
  wire  s_0_179 = m_508_io_s; // @[MUL.scala 262:21]
  wire  c_0_179 = m_508_io_cout; // @[MUL.scala 263:22]
  wire  s_0_180 = m_509_io_s; // @[MUL.scala 262:21]
  wire  c_0_180 = m_509_io_cout; // @[MUL.scala 263:22]
  wire  s_0_181 = m_510_io_s; // @[MUL.scala 262:21]
  wire  c_0_181 = m_510_io_cout; // @[MUL.scala 263:22]
  wire  s_0_182 = m_511_io_s; // @[MUL.scala 262:21]
  wire  c_0_182 = m_511_io_cout; // @[MUL.scala 263:22]
  wire  s_0_183 = m_512_io_s; // @[MUL.scala 262:21]
  wire  c_0_183 = m_512_io_cout; // @[MUL.scala 263:22]
  wire  s_0_184 = m_513_io_s; // @[MUL.scala 262:21]
  wire  c_0_184 = m_513_io_cout; // @[MUL.scala 263:22]
  wire  s_0_185 = m_514_io_s; // @[MUL.scala 262:21]
  wire  c_0_185 = m_514_io_cout; // @[MUL.scala 263:22]
  wire  s_0_186 = m_515_io_s; // @[MUL.scala 262:21]
  wire  c_0_186 = m_515_io_cout; // @[MUL.scala 263:22]
  wire  s_0_187 = m_516_io_s; // @[MUL.scala 262:21]
  wire  c_0_187 = m_516_io_cout; // @[MUL.scala 263:22]
  wire  s_0_188 = m_517_io_s; // @[MUL.scala 262:21]
  wire  c_0_188 = m_517_io_cout; // @[MUL.scala 263:22]
  wire  s_0_189 = m_519_io_s; // @[MUL.scala 262:21]
  wire  c_0_189 = m_519_io_cout; // @[MUL.scala 263:22]
  wire  s_0_190 = m_521_io_s; // @[MUL.scala 262:21]
  wire  c_0_190 = m_521_io_cout; // @[MUL.scala 263:22]
  wire  s_0_191 = m_523_io_s; // @[MUL.scala 262:21]
  wire  c_0_191 = m_523_io_cout; // @[MUL.scala 263:22]
  wire  s_0_192 = m_525_io_s; // @[MUL.scala 262:21]
  wire  c_0_192 = m_525_io_cout; // @[MUL.scala 263:22]
  wire  s_0_193 = m_527_io_s; // @[MUL.scala 262:21]
  wire  c_0_193 = m_527_io_cout; // @[MUL.scala 263:22]
  wire  s_2_122 = m_528_io_s; // @[MUL.scala 262:21]
  wire  c_1_122 = m_528_io_cout; // @[MUL.scala 263:22]
  wire  s_0_194 = m_529_io_s; // @[MUL.scala 262:21]
  wire  c_0_194 = m_529_io_cout; // @[MUL.scala 263:22]
  wire  s_2_123 = m_530_io_s; // @[MUL.scala 262:21]
  wire  c_1_123 = m_530_io_cout; // @[MUL.scala 263:22]
  wire  s_0_195 = m_531_io_s; // @[MUL.scala 262:21]
  wire  c_0_195 = m_531_io_cout; // @[MUL.scala 263:22]
  wire  s_2_124 = m_532_io_s; // @[MUL.scala 262:21]
  wire  c_1_124 = m_532_io_cout; // @[MUL.scala 263:22]
  wire  s_0_196 = m_533_io_s; // @[MUL.scala 262:21]
  wire  c_0_196 = m_533_io_cout; // @[MUL.scala 263:22]
  wire  s_2_125 = m_534_io_s; // @[MUL.scala 262:21]
  wire  c_1_125 = m_534_io_cout; // @[MUL.scala 263:22]
  wire  s_0_197 = m_535_io_s; // @[MUL.scala 262:21]
  wire  c_0_197 = m_535_io_cout; // @[MUL.scala 263:22]
  wire  s_2_126 = m_536_io_s; // @[MUL.scala 262:21]
  wire  c_1_126 = m_536_io_cout; // @[MUL.scala 263:22]
  wire  s_0_198 = m_537_io_s; // @[MUL.scala 262:21]
  wire  c_0_198 = m_537_io_cout; // @[MUL.scala 263:22]
  wire  s_2_127 = m_538_io_s; // @[MUL.scala 262:21]
  wire  c_1_127 = m_538_io_cout; // @[MUL.scala 263:22]
  wire  s_0_199 = m_539_io_s; // @[MUL.scala 262:21]
  wire  c_0_199 = m_539_io_cout; // @[MUL.scala 263:22]
  wire  s_2_128 = m_540_io_s; // @[MUL.scala 262:21]
  wire  c_1_128 = m_540_io_cout; // @[MUL.scala 263:22]
  wire  s_0_200 = m_541_io_s; // @[MUL.scala 262:21]
  wire  c_0_200 = m_541_io_cout; // @[MUL.scala 263:22]
  wire  s_2_129 = m_542_io_s; // @[MUL.scala 262:21]
  wire  c_1_129 = m_542_io_cout; // @[MUL.scala 263:22]
  wire  s_0_201 = m_543_io_s; // @[MUL.scala 262:21]
  wire  c_0_201 = m_543_io_cout; // @[MUL.scala 263:22]
  wire  s_2_130 = m_544_io_s; // @[MUL.scala 262:21]
  wire  c_1_130 = m_544_io_cout; // @[MUL.scala 263:22]
  wire  s_0_202 = m_545_io_s; // @[MUL.scala 262:21]
  wire  c_0_202 = m_545_io_cout; // @[MUL.scala 263:22]
  wire  s_2_131 = m_546_io_s; // @[MUL.scala 262:21]
  wire  c_1_131 = m_546_io_cout; // @[MUL.scala 263:22]
  wire  s_0_203 = m_547_io_s; // @[MUL.scala 262:21]
  wire  c_0_203 = m_547_io_cout; // @[MUL.scala 263:22]
  wire  s_0_204 = m_549_io_s; // @[MUL.scala 262:21]
  wire  c_0_204 = m_549_io_cout; // @[MUL.scala 263:22]
  wire  s_0_205 = m_551_io_s; // @[MUL.scala 262:21]
  wire  c_0_205 = m_551_io_cout; // @[MUL.scala 263:22]
  wire  s_0_206 = m_553_io_s; // @[MUL.scala 262:21]
  wire  c_0_206 = m_553_io_cout; // @[MUL.scala 263:22]
  wire  s_0_207 = m_554_io_s; // @[MUL.scala 262:21]
  wire  c_0_207 = m_554_io_cout; // @[MUL.scala 263:22]
  wire  s_0_208 = m_555_io_s; // @[MUL.scala 262:21]
  wire  c_0_208 = m_555_io_cout; // @[MUL.scala 263:22]
  wire  s_0_209 = m_556_io_s; // @[MUL.scala 262:21]
  wire  c_0_209 = m_556_io_cout; // @[MUL.scala 263:22]
  wire  s_0_210 = m_557_io_s; // @[MUL.scala 262:21]
  wire  c_0_210 = m_557_io_cout; // @[MUL.scala 263:22]
  wire  s_0_211 = m_558_io_s; // @[MUL.scala 262:21]
  wire  c_0_211 = m_558_io_cout; // @[MUL.scala 263:22]
  wire  s_0_212 = m_559_io_s; // @[MUL.scala 262:21]
  wire  c_0_212 = m_559_io_cout; // @[MUL.scala 263:22]
  wire  s_0_213 = m_560_io_s; // @[MUL.scala 262:21]
  wire  c_0_213 = m_560_io_cout; // @[MUL.scala 263:22]
  wire  s_0_214 = m_561_io_s; // @[MUL.scala 262:21]
  wire  c_0_214 = m_561_io_cout; // @[MUL.scala 263:22]
  wire  s_0_215 = m_562_io_s; // @[MUL.scala 262:21]
  wire  c_0_215 = m_562_io_cout; // @[MUL.scala 263:22]
  wire  s_0_216 = m_563_io_s; // @[MUL.scala 262:21]
  wire  c_0_216 = m_563_io_cout; // @[MUL.scala 263:22]
  wire  s_0_217 = m_564_io_s; // @[MUL.scala 262:21]
  wire  c_0_217 = m_564_io_cout; // @[MUL.scala 263:22]
  wire  s_0_218 = m_565_io_s; // @[MUL.scala 262:21]
  wire  c_0_218 = m_565_io_cout; // @[MUL.scala 263:22]
  wire  s_0_219 = m_566_io_s; // @[MUL.scala 262:21]
  wire  c_0_219 = m_566_io_cout; // @[MUL.scala 263:22]
  reg  r_644; // @[Reg.scala 19:16]
  reg  r_645; // @[Reg.scala 19:16]
  reg  r_646; // @[Reg.scala 19:16]
  reg  r_647; // @[Reg.scala 19:16]
  reg  r_648; // @[Reg.scala 19:16]
  reg  r_649; // @[Reg.scala 19:16]
  reg  r_650; // @[Reg.scala 19:16]
  reg  r_651; // @[Reg.scala 19:16]
  reg  r_652; // @[Reg.scala 19:16]
  reg  r_653; // @[Reg.scala 19:16]
  reg  r_654; // @[Reg.scala 19:16]
  reg  r_655; // @[Reg.scala 19:16]
  reg  r_656; // @[Reg.scala 19:16]
  reg  r_657; // @[Reg.scala 19:16]
  reg  r_658; // @[Reg.scala 19:16]
  reg  r_659; // @[Reg.scala 19:16]
  reg  r_660; // @[Reg.scala 19:16]
  reg  r_661; // @[Reg.scala 19:16]
  reg  r_662; // @[Reg.scala 19:16]
  reg  r_663; // @[Reg.scala 19:16]
  reg  r_664; // @[Reg.scala 19:16]
  reg  r_665; // @[Reg.scala 19:16]
  reg  r_666; // @[Reg.scala 19:16]
  reg  r_667; // @[Reg.scala 19:16]
  reg  r_668; // @[Reg.scala 19:16]
  reg  r_669; // @[Reg.scala 19:16]
  reg  r_670; // @[Reg.scala 19:16]
  reg  r_671; // @[Reg.scala 19:16]
  reg  r_672; // @[Reg.scala 19:16]
  reg  r_673; // @[Reg.scala 19:16]
  reg  r_674; // @[Reg.scala 19:16]
  reg  r_675; // @[Reg.scala 19:16]
  reg  r_676; // @[Reg.scala 19:16]
  reg  r_677; // @[Reg.scala 19:16]
  reg  r_678; // @[Reg.scala 19:16]
  reg  r_679; // @[Reg.scala 19:16]
  reg  r_680; // @[Reg.scala 19:16]
  reg  r_681; // @[Reg.scala 19:16]
  reg  r_682; // @[Reg.scala 19:16]
  reg  r_683; // @[Reg.scala 19:16]
  reg  r_684; // @[Reg.scala 19:16]
  reg  r_685; // @[Reg.scala 19:16]
  reg  r_686; // @[Reg.scala 19:16]
  reg  r_687; // @[Reg.scala 19:16]
  reg  r_688; // @[Reg.scala 19:16]
  reg  r_689; // @[Reg.scala 19:16]
  reg  r_690; // @[Reg.scala 19:16]
  reg  r_691; // @[Reg.scala 19:16]
  reg  r_692; // @[Reg.scala 19:16]
  reg  r_693; // @[Reg.scala 19:16]
  reg  r_694; // @[Reg.scala 19:16]
  reg  r_695; // @[Reg.scala 19:16]
  reg  r_696; // @[Reg.scala 19:16]
  reg  r_697; // @[Reg.scala 19:16]
  reg  r_698; // @[Reg.scala 19:16]
  reg  r_699; // @[Reg.scala 19:16]
  reg  r_700; // @[Reg.scala 19:16]
  reg  r_701; // @[Reg.scala 19:16]
  reg  r_702; // @[Reg.scala 19:16]
  reg  r_703; // @[Reg.scala 19:16]
  reg  r_704; // @[Reg.scala 19:16]
  reg  r_705; // @[Reg.scala 19:16]
  reg  r_706; // @[Reg.scala 19:16]
  reg  r_707; // @[Reg.scala 19:16]
  reg  r_708; // @[Reg.scala 19:16]
  reg  r_709; // @[Reg.scala 19:16]
  reg  r_710; // @[Reg.scala 19:16]
  reg  r_711; // @[Reg.scala 19:16]
  reg  r_712; // @[Reg.scala 19:16]
  reg  r_713; // @[Reg.scala 19:16]
  reg  r_714; // @[Reg.scala 19:16]
  reg  r_715; // @[Reg.scala 19:16]
  reg  r_716; // @[Reg.scala 19:16]
  reg  r_717; // @[Reg.scala 19:16]
  reg  r_718; // @[Reg.scala 19:16]
  reg  r_719; // @[Reg.scala 19:16]
  reg  r_720; // @[Reg.scala 19:16]
  reg  r_721; // @[Reg.scala 19:16]
  reg  r_722; // @[Reg.scala 19:16]
  reg  r_723; // @[Reg.scala 19:16]
  reg  r_724; // @[Reg.scala 19:16]
  reg  r_725; // @[Reg.scala 19:16]
  reg  r_726; // @[Reg.scala 19:16]
  reg  r_727; // @[Reg.scala 19:16]
  reg  r_728; // @[Reg.scala 19:16]
  reg  r_729; // @[Reg.scala 19:16]
  reg  r_730; // @[Reg.scala 19:16]
  reg  r_731; // @[Reg.scala 19:16]
  reg  r_732; // @[Reg.scala 19:16]
  reg  r_733; // @[Reg.scala 19:16]
  reg  r_734; // @[Reg.scala 19:16]
  reg  r_735; // @[Reg.scala 19:16]
  reg  r_736; // @[Reg.scala 19:16]
  reg  r_737; // @[Reg.scala 19:16]
  reg  r_738; // @[Reg.scala 19:16]
  reg  r_739; // @[Reg.scala 19:16]
  reg  r_740; // @[Reg.scala 19:16]
  reg  r_741; // @[Reg.scala 19:16]
  reg  r_742; // @[Reg.scala 19:16]
  reg  r_743; // @[Reg.scala 19:16]
  reg  r_744; // @[Reg.scala 19:16]
  reg  r_745; // @[Reg.scala 19:16]
  reg  r_746; // @[Reg.scala 19:16]
  reg  r_747; // @[Reg.scala 19:16]
  reg  r_748; // @[Reg.scala 19:16]
  reg  r_749; // @[Reg.scala 19:16]
  reg  r_750; // @[Reg.scala 19:16]
  reg  r_751; // @[Reg.scala 19:16]
  reg  r_752; // @[Reg.scala 19:16]
  reg  r_753; // @[Reg.scala 19:16]
  reg  r_754; // @[Reg.scala 19:16]
  reg  r_755; // @[Reg.scala 19:16]
  reg  r_756; // @[Reg.scala 19:16]
  reg  r_757; // @[Reg.scala 19:16]
  reg  r_758; // @[Reg.scala 19:16]
  reg  r_759; // @[Reg.scala 19:16]
  reg  r_760; // @[Reg.scala 19:16]
  reg  r_761; // @[Reg.scala 19:16]
  reg  r_762; // @[Reg.scala 19:16]
  reg  r_763; // @[Reg.scala 19:16]
  reg  r_764; // @[Reg.scala 19:16]
  reg  r_765; // @[Reg.scala 19:16]
  reg  r_766; // @[Reg.scala 19:16]
  reg  r_767; // @[Reg.scala 19:16]
  reg  r_768; // @[Reg.scala 19:16]
  reg  r_769; // @[Reg.scala 19:16]
  reg  r_770; // @[Reg.scala 19:16]
  reg  r_771; // @[Reg.scala 19:16]
  reg  r_772; // @[Reg.scala 19:16]
  reg  r_773; // @[Reg.scala 19:16]
  reg  r_774; // @[Reg.scala 19:16]
  reg  r_775; // @[Reg.scala 19:16]
  reg  r_776; // @[Reg.scala 19:16]
  reg  r_777; // @[Reg.scala 19:16]
  reg  r_778; // @[Reg.scala 19:16]
  reg  r_779; // @[Reg.scala 19:16]
  reg  r_780; // @[Reg.scala 19:16]
  reg  r_781; // @[Reg.scala 19:16]
  reg  r_782; // @[Reg.scala 19:16]
  reg  r_783; // @[Reg.scala 19:16]
  reg  r_784; // @[Reg.scala 19:16]
  reg  r_785; // @[Reg.scala 19:16]
  reg  r_786; // @[Reg.scala 19:16]
  reg  r_787; // @[Reg.scala 19:16]
  reg  r_788; // @[Reg.scala 19:16]
  reg  r_789; // @[Reg.scala 19:16]
  reg  r_790; // @[Reg.scala 19:16]
  reg  r_791; // @[Reg.scala 19:16]
  reg  r_792; // @[Reg.scala 19:16]
  reg  r_793; // @[Reg.scala 19:16]
  reg  r_794; // @[Reg.scala 19:16]
  reg  r_795; // @[Reg.scala 19:16]
  reg  r_796; // @[Reg.scala 19:16]
  reg  r_797; // @[Reg.scala 19:16]
  reg  r_798; // @[Reg.scala 19:16]
  reg  r_799; // @[Reg.scala 19:16]
  reg  r_800; // @[Reg.scala 19:16]
  reg  r_801; // @[Reg.scala 19:16]
  reg  r_802; // @[Reg.scala 19:16]
  reg  r_803; // @[Reg.scala 19:16]
  reg  r_804; // @[Reg.scala 19:16]
  reg  r_805; // @[Reg.scala 19:16]
  reg  r_806; // @[Reg.scala 19:16]
  reg  r_807; // @[Reg.scala 19:16]
  reg  r_808; // @[Reg.scala 19:16]
  reg  r_809; // @[Reg.scala 19:16]
  reg  r_810; // @[Reg.scala 19:16]
  reg  r_811; // @[Reg.scala 19:16]
  reg  r_812; // @[Reg.scala 19:16]
  reg  r_813; // @[Reg.scala 19:16]
  reg  r_814; // @[Reg.scala 19:16]
  reg  r_815; // @[Reg.scala 19:16]
  reg  r_816; // @[Reg.scala 19:16]
  reg  r_817; // @[Reg.scala 19:16]
  reg  r_818; // @[Reg.scala 19:16]
  reg  r_819; // @[Reg.scala 19:16]
  reg  r_820; // @[Reg.scala 19:16]
  reg  r_821; // @[Reg.scala 19:16]
  reg  r_822; // @[Reg.scala 19:16]
  reg  r_823; // @[Reg.scala 19:16]
  reg  r_824; // @[Reg.scala 19:16]
  reg  r_825; // @[Reg.scala 19:16]
  wire  s_0_254 = m_661_io_s; // @[MUL.scala 262:21]
  wire  c_0_254 = m_661_io_cout; // @[MUL.scala 263:22]
  wire  s_0_255 = m_662_io_s; // @[MUL.scala 262:21]
  wire  c_0_255 = m_662_io_cout; // @[MUL.scala 263:22]
  wire  s_0_256 = m_663_io_s; // @[MUL.scala 262:21]
  wire  c_0_256 = m_663_io_cout; // @[MUL.scala 263:22]
  wire  s_0_257 = m_664_io_s; // @[MUL.scala 262:21]
  wire  c_0_257 = m_664_io_cout; // @[MUL.scala 263:22]
  wire  s_0_258 = m_665_io_s; // @[MUL.scala 262:21]
  wire  c_0_258 = m_665_io_cout; // @[MUL.scala 263:22]
  wire  s_0_259 = m_666_io_s; // @[MUL.scala 262:21]
  wire  c_0_259 = m_666_io_cout; // @[MUL.scala 263:22]
  wire  s_0_260 = m_667_io_s; // @[MUL.scala 262:21]
  wire  c_0_260 = m_667_io_cout; // @[MUL.scala 263:22]
  wire  s_0_261 = m_668_io_s; // @[MUL.scala 262:21]
  wire  c_0_261 = m_668_io_cout; // @[MUL.scala 263:22]
  wire  s_0_262 = m_669_io_s; // @[MUL.scala 262:21]
  wire  c_0_262 = m_669_io_cout; // @[MUL.scala 263:22]
  wire  s_0_263 = m_670_io_s; // @[MUL.scala 262:21]
  wire  c_0_263 = m_670_io_cout; // @[MUL.scala 263:22]
  wire  s_0_264 = m_671_io_s; // @[MUL.scala 262:21]
  wire  c_0_264 = m_671_io_cout; // @[MUL.scala 263:22]
  wire  s_0_265 = m_672_io_s; // @[MUL.scala 262:21]
  wire  c_0_265 = m_672_io_cout; // @[MUL.scala 263:22]
  wire  s_0_266 = m_673_io_s; // @[MUL.scala 262:21]
  wire  c_0_266 = m_673_io_cout; // @[MUL.scala 263:22]
  wire  s_0_267 = m_674_io_s; // @[MUL.scala 262:21]
  wire  c_0_267 = m_674_io_cout; // @[MUL.scala 263:22]
  wire  s_0_268 = m_675_io_s; // @[MUL.scala 262:21]
  wire  c_0_268 = m_675_io_cout; // @[MUL.scala 263:22]
  wire  s_0_269 = m_676_io_s; // @[MUL.scala 262:21]
  wire  c_0_269 = m_676_io_cout; // @[MUL.scala 263:22]
  wire  s_0_270 = m_677_io_s; // @[MUL.scala 262:21]
  wire  c_0_270 = m_677_io_cout; // @[MUL.scala 263:22]
  wire  s_0_271 = m_678_io_s; // @[MUL.scala 262:21]
  wire  c_0_271 = m_678_io_cout; // @[MUL.scala 263:22]
  wire [7:0] sum_lo_lo_lo = {m_642_io_out_0,m_641_io_out_0,m_640_io_out_0,m_577_io_out_0,r_647,r_646,r_645,r_644}; // @[Cat.scala 33:92]
  wire [7:0] sum_lo_hi_lo = {m_658_io_out_0,m_657_io_out_0,m_656_io_out_0,m_655_io_out_0,m_654_io_out_0,m_653_io_out_0,
    m_652_io_out_0,m_651_io_out_0}; // @[Cat.scala 33:92]
  wire [16:0] sum_lo_hi = {s_0_260,s_0_259,s_0_258,s_0_257,s_0_256,s_0_255,s_0_254,m_660_io_out_0,m_659_io_out_0,
    sum_lo_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] sum_lo = {sum_lo_hi,m_650_io_out_0,m_649_io_out_0,m_648_io_out_0,m_647_io_out_0,m_646_io_out_0,
    m_645_io_out_0,m_644_io_out_0,m_643_io_out_0,sum_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] sum_hi_lo_lo = {s_0_268,s_0_267,s_0_266,s_0_265,s_0_264,s_0_263,s_0_262,s_0_261}; // @[Cat.scala 33:92]
  wire [16:0] sum_hi_lo = {m_684_io_out_0,m_683_io_out_0,m_682_io_out_0,m_681_io_out_0,m_680_io_out_0,m_679_io_out_0,
    s_0_271,s_0_270,s_0_269,sum_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] sum_hi_hi_lo = {m_692_io_out_0,m_691_io_out_0,m_690_io_out_0,m_689_io_out_0,m_688_io_out_0,m_687_io_out_0,
    m_686_io_out_0,m_685_io_out_0}; // @[Cat.scala 33:92]
  wire [16:0] sum_hi_hi = {m_701_io_out_0,m_700_io_out_0,m_699_io_out_0,m_698_io_out_0,m_697_io_out_0,m_696_io_out_0,
    m_695_io_out_0,m_694_io_out_0,m_693_io_out_0,sum_hi_hi_lo}; // @[Cat.scala 33:92]
  wire [66:0] sum = {sum_hi_hi,sum_hi_lo,sum_lo}; // @[Cat.scala 33:92]
  wire [6:0] carry_lo_lo_lo = {m_646_io_out_1,m_645_io_out_1,m_644_io_out_1,m_643_io_out_1,m_642_io_out_1,m_641_io_out_1
    ,m_640_io_out_1}; // @[Cat.scala 33:92]
  wire [14:0] carry_lo_lo = {m_654_io_out_1,m_653_io_out_1,m_652_io_out_1,m_651_io_out_1,m_650_io_out_1,m_649_io_out_1,
    m_648_io_out_1,m_647_io_out_1,carry_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [6:0] carry_lo_hi_lo = {c_0_254,m_660_io_out_1,m_659_io_out_1,m_658_io_out_1,m_657_io_out_1,m_656_io_out_1,
    m_655_io_out_1}; // @[Cat.scala 33:92]
  wire [29:0] carry_lo = {c_0_262,c_0_261,c_0_260,c_0_259,c_0_258,c_0_257,c_0_256,c_0_255,carry_lo_hi_lo,carry_lo_lo}; // @[Cat.scala 33:92]
  wire [6:0] carry_hi_lo_lo = {c_0_269,c_0_268,c_0_267,c_0_266,c_0_265,c_0_264,c_0_263}; // @[Cat.scala 33:92]
  wire [14:0] carry_hi_lo = {m_684_io_out_1,m_683_io_out_1,m_682_io_out_1,m_681_io_out_1,m_680_io_out_1,m_679_io_out_1,
    c_0_271,c_0_270,carry_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] carry_hi_hi_lo = {m_692_io_out_1,m_691_io_out_1,m_690_io_out_1,m_689_io_out_1,m_688_io_out_1,m_687_io_out_1
    ,m_686_io_out_1,m_685_io_out_1}; // @[Cat.scala 33:92]
  wire [30:0] carry_hi = {m_700_io_out_1,m_699_io_out_1,m_698_io_out_1,m_697_io_out_1,m_696_io_out_1,m_695_io_out_1,
    m_694_io_out_1,m_693_io_out_1,carry_hi_hi_lo,carry_hi_lo}; // @[Cat.scala 33:92]
  wire [66:0] cout = {carry_hi,carry_lo,6'h0}; // @[Cat.scala 33:92]
  wire [66:0] result = sum + cout; // @[MUL.scala 342:20]
  reg [7:0] count; // @[MUL.scala 344:22]
  wire [7:0] _count_T_5 = count + 8'h1; // @[MUL.scala 346:81]
  Improved_Partial_product m ( // @[MUL.scala 81:21]
    .io_y_3(m_io_y_3),
    .io_x(m_io_x),
    .io_p(m_io_p),
    .io_carry(m_io_carry)
  );
  Improved_Partial_product m_1 ( // @[MUL.scala 81:21]
    .io_y_3(m_1_io_y_3),
    .io_x(m_1_io_x),
    .io_p(m_1_io_p),
    .io_carry(m_1_io_carry)
  );
  Improved_Partial_product m_2 ( // @[MUL.scala 81:21]
    .io_y_3(m_2_io_y_3),
    .io_x(m_2_io_x),
    .io_p(m_2_io_p),
    .io_carry(m_2_io_carry)
  );
  Improved_Partial_product m_3 ( // @[MUL.scala 81:21]
    .io_y_3(m_3_io_y_3),
    .io_x(m_3_io_x),
    .io_p(m_3_io_p),
    .io_carry(m_3_io_carry)
  );
  Improved_Partial_product m_4 ( // @[MUL.scala 81:21]
    .io_y_3(m_4_io_y_3),
    .io_x(m_4_io_x),
    .io_p(m_4_io_p),
    .io_carry(m_4_io_carry)
  );
  Improved_Partial_product m_5 ( // @[MUL.scala 81:21]
    .io_y_3(m_5_io_y_3),
    .io_x(m_5_io_x),
    .io_p(m_5_io_p),
    .io_carry(m_5_io_carry)
  );
  Improved_Partial_product m_6 ( // @[MUL.scala 81:21]
    .io_y_3(m_6_io_y_3),
    .io_x(m_6_io_x),
    .io_p(m_6_io_p),
    .io_carry(m_6_io_carry)
  );
  Improved_Partial_product m_7 ( // @[MUL.scala 81:21]
    .io_y_3(m_7_io_y_3),
    .io_x(m_7_io_x),
    .io_p(m_7_io_p),
    .io_carry(m_7_io_carry)
  );
  Improved_Partial_product m_8 ( // @[MUL.scala 81:21]
    .io_y_3(m_8_io_y_3),
    .io_x(m_8_io_x),
    .io_p(m_8_io_p),
    .io_carry(m_8_io_carry)
  );
  Improved_Partial_product m_9 ( // @[MUL.scala 81:21]
    .io_y_3(m_9_io_y_3),
    .io_x(m_9_io_x),
    .io_p(m_9_io_p),
    .io_carry(m_9_io_carry)
  );
  Improved_Partial_product m_10 ( // @[MUL.scala 81:21]
    .io_y_3(m_10_io_y_3),
    .io_x(m_10_io_x),
    .io_p(m_10_io_p),
    .io_carry(m_10_io_carry)
  );
  Improved_Partial_product m_11 ( // @[MUL.scala 81:21]
    .io_y_3(m_11_io_y_3),
    .io_x(m_11_io_x),
    .io_p(m_11_io_p),
    .io_carry(m_11_io_carry)
  );
  Improved_Partial_product m_12 ( // @[MUL.scala 81:21]
    .io_y_3(m_12_io_y_3),
    .io_x(m_12_io_x),
    .io_p(m_12_io_p),
    .io_carry(m_12_io_carry)
  );
  Improved_Partial_product m_13 ( // @[MUL.scala 81:21]
    .io_y_3(m_13_io_y_3),
    .io_x(m_13_io_x),
    .io_p(m_13_io_p),
    .io_carry(m_13_io_carry)
  );
  Improved_Partial_product m_14 ( // @[MUL.scala 81:21]
    .io_y_3(m_14_io_y_3),
    .io_x(m_14_io_x),
    .io_p(m_14_io_p),
    .io_carry(m_14_io_carry)
  );
  Improved_Partial_product m_15 ( // @[MUL.scala 81:21]
    .io_y_3(m_15_io_y_3),
    .io_x(m_15_io_x),
    .io_p(m_15_io_p),
    .io_carry(m_15_io_carry)
  );
  Improved_Partial_product m_16 ( // @[MUL.scala 81:21]
    .io_y_3(m_16_io_y_3),
    .io_x(m_16_io_x),
    .io_p(m_16_io_p),
    .io_carry(m_16_io_carry)
  );
  Half_Adder m_17 ( // @[MUL.scala 124:19]
    .io_in_0(m_17_io_in_0),
    .io_in_1(m_17_io_in_1),
    .io_out_0(m_17_io_out_0),
    .io_out_1(m_17_io_out_1)
  );
  Half_Adder m_18 ( // @[MUL.scala 124:19]
    .io_in_0(m_18_io_in_0),
    .io_in_1(m_18_io_in_1),
    .io_out_0(m_18_io_out_0),
    .io_out_1(m_18_io_out_1)
  );
  Adder m_19 ( // @[MUL.scala 102:19]
    .io_x1(m_19_io_x1),
    .io_x2(m_19_io_x2),
    .io_x3(m_19_io_x3),
    .io_s(m_19_io_s),
    .io_cout(m_19_io_cout)
  );
  Adder m_20 ( // @[MUL.scala 102:19]
    .io_x1(m_20_io_x1),
    .io_x2(m_20_io_x2),
    .io_x3(m_20_io_x3),
    .io_s(m_20_io_s),
    .io_cout(m_20_io_cout)
  );
  Adder m_21 ( // @[MUL.scala 102:19]
    .io_x1(m_21_io_x1),
    .io_x2(m_21_io_x2),
    .io_x3(m_21_io_x3),
    .io_s(m_21_io_s),
    .io_cout(m_21_io_cout)
  );
  Adder m_22 ( // @[MUL.scala 102:19]
    .io_x1(m_22_io_x1),
    .io_x2(m_22_io_x2),
    .io_x3(m_22_io_x3),
    .io_s(m_22_io_s),
    .io_cout(m_22_io_cout)
  );
  Adder m_23 ( // @[MUL.scala 102:19]
    .io_x1(m_23_io_x1),
    .io_x2(m_23_io_x2),
    .io_x3(m_23_io_x3),
    .io_s(m_23_io_s),
    .io_cout(m_23_io_cout)
  );
  Half_Adder m_24 ( // @[MUL.scala 124:19]
    .io_in_0(m_24_io_in_0),
    .io_in_1(m_24_io_in_1),
    .io_out_0(m_24_io_out_0),
    .io_out_1(m_24_io_out_1)
  );
  Adder m_25 ( // @[MUL.scala 102:19]
    .io_x1(m_25_io_x1),
    .io_x2(m_25_io_x2),
    .io_x3(m_25_io_x3),
    .io_s(m_25_io_s),
    .io_cout(m_25_io_cout)
  );
  Half_Adder m_26 ( // @[MUL.scala 124:19]
    .io_in_0(m_26_io_in_0),
    .io_in_1(m_26_io_in_1),
    .io_out_0(m_26_io_out_0),
    .io_out_1(m_26_io_out_1)
  );
  Adder m_27 ( // @[MUL.scala 102:19]
    .io_x1(m_27_io_x1),
    .io_x2(m_27_io_x2),
    .io_x3(m_27_io_x3),
    .io_s(m_27_io_s),
    .io_cout(m_27_io_cout)
  );
  Adder m_28 ( // @[MUL.scala 102:19]
    .io_x1(m_28_io_x1),
    .io_x2(m_28_io_x2),
    .io_x3(m_28_io_x3),
    .io_s(m_28_io_s),
    .io_cout(m_28_io_cout)
  );
  Adder m_29 ( // @[MUL.scala 102:19]
    .io_x1(m_29_io_x1),
    .io_x2(m_29_io_x2),
    .io_x3(m_29_io_x3),
    .io_s(m_29_io_s),
    .io_cout(m_29_io_cout)
  );
  Adder m_30 ( // @[MUL.scala 102:19]
    .io_x1(m_30_io_x1),
    .io_x2(m_30_io_x2),
    .io_x3(m_30_io_x3),
    .io_s(m_30_io_s),
    .io_cout(m_30_io_cout)
  );
  Adder m_31 ( // @[MUL.scala 102:19]
    .io_x1(m_31_io_x1),
    .io_x2(m_31_io_x2),
    .io_x3(m_31_io_x3),
    .io_s(m_31_io_s),
    .io_cout(m_31_io_cout)
  );
  Adder m_32 ( // @[MUL.scala 102:19]
    .io_x1(m_32_io_x1),
    .io_x2(m_32_io_x2),
    .io_x3(m_32_io_x3),
    .io_s(m_32_io_s),
    .io_cout(m_32_io_cout)
  );
  Adder m_33 ( // @[MUL.scala 102:19]
    .io_x1(m_33_io_x1),
    .io_x2(m_33_io_x2),
    .io_x3(m_33_io_x3),
    .io_s(m_33_io_s),
    .io_cout(m_33_io_cout)
  );
  Adder m_34 ( // @[MUL.scala 102:19]
    .io_x1(m_34_io_x1),
    .io_x2(m_34_io_x2),
    .io_x3(m_34_io_x3),
    .io_s(m_34_io_s),
    .io_cout(m_34_io_cout)
  );
  Adder m_35 ( // @[MUL.scala 102:19]
    .io_x1(m_35_io_x1),
    .io_x2(m_35_io_x2),
    .io_x3(m_35_io_x3),
    .io_s(m_35_io_s),
    .io_cout(m_35_io_cout)
  );
  Adder m_36 ( // @[MUL.scala 102:19]
    .io_x1(m_36_io_x1),
    .io_x2(m_36_io_x2),
    .io_x3(m_36_io_x3),
    .io_s(m_36_io_s),
    .io_cout(m_36_io_cout)
  );
  Half_Adder m_37 ( // @[MUL.scala 124:19]
    .io_in_0(m_37_io_in_0),
    .io_in_1(m_37_io_in_1),
    .io_out_0(m_37_io_out_0),
    .io_out_1(m_37_io_out_1)
  );
  Adder m_38 ( // @[MUL.scala 102:19]
    .io_x1(m_38_io_x1),
    .io_x2(m_38_io_x2),
    .io_x3(m_38_io_x3),
    .io_s(m_38_io_s),
    .io_cout(m_38_io_cout)
  );
  Adder m_39 ( // @[MUL.scala 102:19]
    .io_x1(m_39_io_x1),
    .io_x2(m_39_io_x2),
    .io_x3(m_39_io_x3),
    .io_s(m_39_io_s),
    .io_cout(m_39_io_cout)
  );
  Half_Adder m_40 ( // @[MUL.scala 124:19]
    .io_in_0(m_40_io_in_0),
    .io_in_1(m_40_io_in_1),
    .io_out_0(m_40_io_out_0),
    .io_out_1(m_40_io_out_1)
  );
  Adder m_41 ( // @[MUL.scala 102:19]
    .io_x1(m_41_io_x1),
    .io_x2(m_41_io_x2),
    .io_x3(m_41_io_x3),
    .io_s(m_41_io_s),
    .io_cout(m_41_io_cout)
  );
  Adder m_42 ( // @[MUL.scala 102:19]
    .io_x1(m_42_io_x1),
    .io_x2(m_42_io_x2),
    .io_x3(m_42_io_x3),
    .io_s(m_42_io_s),
    .io_cout(m_42_io_cout)
  );
  Adder m_43 ( // @[MUL.scala 102:19]
    .io_x1(m_43_io_x1),
    .io_x2(m_43_io_x2),
    .io_x3(m_43_io_x3),
    .io_s(m_43_io_s),
    .io_cout(m_43_io_cout)
  );
  Adder m_44 ( // @[MUL.scala 102:19]
    .io_x1(m_44_io_x1),
    .io_x2(m_44_io_x2),
    .io_x3(m_44_io_x3),
    .io_s(m_44_io_s),
    .io_cout(m_44_io_cout)
  );
  Adder m_45 ( // @[MUL.scala 102:19]
    .io_x1(m_45_io_x1),
    .io_x2(m_45_io_x2),
    .io_x3(m_45_io_x3),
    .io_s(m_45_io_s),
    .io_cout(m_45_io_cout)
  );
  Adder m_46 ( // @[MUL.scala 102:19]
    .io_x1(m_46_io_x1),
    .io_x2(m_46_io_x2),
    .io_x3(m_46_io_x3),
    .io_s(m_46_io_s),
    .io_cout(m_46_io_cout)
  );
  Adder m_47 ( // @[MUL.scala 102:19]
    .io_x1(m_47_io_x1),
    .io_x2(m_47_io_x2),
    .io_x3(m_47_io_x3),
    .io_s(m_47_io_s),
    .io_cout(m_47_io_cout)
  );
  Adder m_48 ( // @[MUL.scala 102:19]
    .io_x1(m_48_io_x1),
    .io_x2(m_48_io_x2),
    .io_x3(m_48_io_x3),
    .io_s(m_48_io_s),
    .io_cout(m_48_io_cout)
  );
  Adder m_49 ( // @[MUL.scala 102:19]
    .io_x1(m_49_io_x1),
    .io_x2(m_49_io_x2),
    .io_x3(m_49_io_x3),
    .io_s(m_49_io_s),
    .io_cout(m_49_io_cout)
  );
  Adder m_50 ( // @[MUL.scala 102:19]
    .io_x1(m_50_io_x1),
    .io_x2(m_50_io_x2),
    .io_x3(m_50_io_x3),
    .io_s(m_50_io_s),
    .io_cout(m_50_io_cout)
  );
  Adder m_51 ( // @[MUL.scala 102:19]
    .io_x1(m_51_io_x1),
    .io_x2(m_51_io_x2),
    .io_x3(m_51_io_x3),
    .io_s(m_51_io_s),
    .io_cout(m_51_io_cout)
  );
  Adder m_52 ( // @[MUL.scala 102:19]
    .io_x1(m_52_io_x1),
    .io_x2(m_52_io_x2),
    .io_x3(m_52_io_x3),
    .io_s(m_52_io_s),
    .io_cout(m_52_io_cout)
  );
  Adder m_53 ( // @[MUL.scala 102:19]
    .io_x1(m_53_io_x1),
    .io_x2(m_53_io_x2),
    .io_x3(m_53_io_x3),
    .io_s(m_53_io_s),
    .io_cout(m_53_io_cout)
  );
  Adder m_54 ( // @[MUL.scala 102:19]
    .io_x1(m_54_io_x1),
    .io_x2(m_54_io_x2),
    .io_x3(m_54_io_x3),
    .io_s(m_54_io_s),
    .io_cout(m_54_io_cout)
  );
  Adder m_55 ( // @[MUL.scala 102:19]
    .io_x1(m_55_io_x1),
    .io_x2(m_55_io_x2),
    .io_x3(m_55_io_x3),
    .io_s(m_55_io_s),
    .io_cout(m_55_io_cout)
  );
  Half_Adder m_56 ( // @[MUL.scala 124:19]
    .io_in_0(m_56_io_in_0),
    .io_in_1(m_56_io_in_1),
    .io_out_0(m_56_io_out_0),
    .io_out_1(m_56_io_out_1)
  );
  Adder m_57 ( // @[MUL.scala 102:19]
    .io_x1(m_57_io_x1),
    .io_x2(m_57_io_x2),
    .io_x3(m_57_io_x3),
    .io_s(m_57_io_s),
    .io_cout(m_57_io_cout)
  );
  Adder m_58 ( // @[MUL.scala 102:19]
    .io_x1(m_58_io_x1),
    .io_x2(m_58_io_x2),
    .io_x3(m_58_io_x3),
    .io_s(m_58_io_s),
    .io_cout(m_58_io_cout)
  );
  Adder m_59 ( // @[MUL.scala 102:19]
    .io_x1(m_59_io_x1),
    .io_x2(m_59_io_x2),
    .io_x3(m_59_io_x3),
    .io_s(m_59_io_s),
    .io_cout(m_59_io_cout)
  );
  Half_Adder m_60 ( // @[MUL.scala 124:19]
    .io_in_0(m_60_io_in_0),
    .io_in_1(m_60_io_in_1),
    .io_out_0(m_60_io_out_0),
    .io_out_1(m_60_io_out_1)
  );
  Adder m_61 ( // @[MUL.scala 102:19]
    .io_x1(m_61_io_x1),
    .io_x2(m_61_io_x2),
    .io_x3(m_61_io_x3),
    .io_s(m_61_io_s),
    .io_cout(m_61_io_cout)
  );
  Adder m_62 ( // @[MUL.scala 102:19]
    .io_x1(m_62_io_x1),
    .io_x2(m_62_io_x2),
    .io_x3(m_62_io_x3),
    .io_s(m_62_io_s),
    .io_cout(m_62_io_cout)
  );
  Adder m_63 ( // @[MUL.scala 102:19]
    .io_x1(m_63_io_x1),
    .io_x2(m_63_io_x2),
    .io_x3(m_63_io_x3),
    .io_s(m_63_io_s),
    .io_cout(m_63_io_cout)
  );
  Adder m_64 ( // @[MUL.scala 102:19]
    .io_x1(m_64_io_x1),
    .io_x2(m_64_io_x2),
    .io_x3(m_64_io_x3),
    .io_s(m_64_io_s),
    .io_cout(m_64_io_cout)
  );
  Adder m_65 ( // @[MUL.scala 102:19]
    .io_x1(m_65_io_x1),
    .io_x2(m_65_io_x2),
    .io_x3(m_65_io_x3),
    .io_s(m_65_io_s),
    .io_cout(m_65_io_cout)
  );
  Adder m_66 ( // @[MUL.scala 102:19]
    .io_x1(m_66_io_x1),
    .io_x2(m_66_io_x2),
    .io_x3(m_66_io_x3),
    .io_s(m_66_io_s),
    .io_cout(m_66_io_cout)
  );
  Adder m_67 ( // @[MUL.scala 102:19]
    .io_x1(m_67_io_x1),
    .io_x2(m_67_io_x2),
    .io_x3(m_67_io_x3),
    .io_s(m_67_io_s),
    .io_cout(m_67_io_cout)
  );
  Adder m_68 ( // @[MUL.scala 102:19]
    .io_x1(m_68_io_x1),
    .io_x2(m_68_io_x2),
    .io_x3(m_68_io_x3),
    .io_s(m_68_io_s),
    .io_cout(m_68_io_cout)
  );
  Adder m_69 ( // @[MUL.scala 102:19]
    .io_x1(m_69_io_x1),
    .io_x2(m_69_io_x2),
    .io_x3(m_69_io_x3),
    .io_s(m_69_io_s),
    .io_cout(m_69_io_cout)
  );
  Adder m_70 ( // @[MUL.scala 102:19]
    .io_x1(m_70_io_x1),
    .io_x2(m_70_io_x2),
    .io_x3(m_70_io_x3),
    .io_s(m_70_io_s),
    .io_cout(m_70_io_cout)
  );
  Adder m_71 ( // @[MUL.scala 102:19]
    .io_x1(m_71_io_x1),
    .io_x2(m_71_io_x2),
    .io_x3(m_71_io_x3),
    .io_s(m_71_io_s),
    .io_cout(m_71_io_cout)
  );
  Adder m_72 ( // @[MUL.scala 102:19]
    .io_x1(m_72_io_x1),
    .io_x2(m_72_io_x2),
    .io_x3(m_72_io_x3),
    .io_s(m_72_io_s),
    .io_cout(m_72_io_cout)
  );
  Adder m_73 ( // @[MUL.scala 102:19]
    .io_x1(m_73_io_x1),
    .io_x2(m_73_io_x2),
    .io_x3(m_73_io_x3),
    .io_s(m_73_io_s),
    .io_cout(m_73_io_cout)
  );
  Adder m_74 ( // @[MUL.scala 102:19]
    .io_x1(m_74_io_x1),
    .io_x2(m_74_io_x2),
    .io_x3(m_74_io_x3),
    .io_s(m_74_io_s),
    .io_cout(m_74_io_cout)
  );
  Adder m_75 ( // @[MUL.scala 102:19]
    .io_x1(m_75_io_x1),
    .io_x2(m_75_io_x2),
    .io_x3(m_75_io_x3),
    .io_s(m_75_io_s),
    .io_cout(m_75_io_cout)
  );
  Adder m_76 ( // @[MUL.scala 102:19]
    .io_x1(m_76_io_x1),
    .io_x2(m_76_io_x2),
    .io_x3(m_76_io_x3),
    .io_s(m_76_io_s),
    .io_cout(m_76_io_cout)
  );
  Adder m_77 ( // @[MUL.scala 102:19]
    .io_x1(m_77_io_x1),
    .io_x2(m_77_io_x2),
    .io_x3(m_77_io_x3),
    .io_s(m_77_io_s),
    .io_cout(m_77_io_cout)
  );
  Adder m_78 ( // @[MUL.scala 102:19]
    .io_x1(m_78_io_x1),
    .io_x2(m_78_io_x2),
    .io_x3(m_78_io_x3),
    .io_s(m_78_io_s),
    .io_cout(m_78_io_cout)
  );
  Adder m_79 ( // @[MUL.scala 102:19]
    .io_x1(m_79_io_x1),
    .io_x2(m_79_io_x2),
    .io_x3(m_79_io_x3),
    .io_s(m_79_io_s),
    .io_cout(m_79_io_cout)
  );
  Adder m_80 ( // @[MUL.scala 102:19]
    .io_x1(m_80_io_x1),
    .io_x2(m_80_io_x2),
    .io_x3(m_80_io_x3),
    .io_s(m_80_io_s),
    .io_cout(m_80_io_cout)
  );
  Half_Adder m_81 ( // @[MUL.scala 124:19]
    .io_in_0(m_81_io_in_0),
    .io_in_1(m_81_io_in_1),
    .io_out_0(m_81_io_out_0),
    .io_out_1(m_81_io_out_1)
  );
  Adder m_82 ( // @[MUL.scala 102:19]
    .io_x1(m_82_io_x1),
    .io_x2(m_82_io_x2),
    .io_x3(m_82_io_x3),
    .io_s(m_82_io_s),
    .io_cout(m_82_io_cout)
  );
  Adder m_83 ( // @[MUL.scala 102:19]
    .io_x1(m_83_io_x1),
    .io_x2(m_83_io_x2),
    .io_x3(m_83_io_x3),
    .io_s(m_83_io_s),
    .io_cout(m_83_io_cout)
  );
  Adder m_84 ( // @[MUL.scala 102:19]
    .io_x1(m_84_io_x1),
    .io_x2(m_84_io_x2),
    .io_x3(m_84_io_x3),
    .io_s(m_84_io_s),
    .io_cout(m_84_io_cout)
  );
  Adder m_85 ( // @[MUL.scala 102:19]
    .io_x1(m_85_io_x1),
    .io_x2(m_85_io_x2),
    .io_x3(m_85_io_x3),
    .io_s(m_85_io_s),
    .io_cout(m_85_io_cout)
  );
  Half_Adder m_86 ( // @[MUL.scala 124:19]
    .io_in_0(m_86_io_in_0),
    .io_in_1(m_86_io_in_1),
    .io_out_0(m_86_io_out_0),
    .io_out_1(m_86_io_out_1)
  );
  Adder m_87 ( // @[MUL.scala 102:19]
    .io_x1(m_87_io_x1),
    .io_x2(m_87_io_x2),
    .io_x3(m_87_io_x3),
    .io_s(m_87_io_s),
    .io_cout(m_87_io_cout)
  );
  Adder m_88 ( // @[MUL.scala 102:19]
    .io_x1(m_88_io_x1),
    .io_x2(m_88_io_x2),
    .io_x3(m_88_io_x3),
    .io_s(m_88_io_s),
    .io_cout(m_88_io_cout)
  );
  Adder m_89 ( // @[MUL.scala 102:19]
    .io_x1(m_89_io_x1),
    .io_x2(m_89_io_x2),
    .io_x3(m_89_io_x3),
    .io_s(m_89_io_s),
    .io_cout(m_89_io_cout)
  );
  Adder m_90 ( // @[MUL.scala 102:19]
    .io_x1(m_90_io_x1),
    .io_x2(m_90_io_x2),
    .io_x3(m_90_io_x3),
    .io_s(m_90_io_s),
    .io_cout(m_90_io_cout)
  );
  Adder m_91 ( // @[MUL.scala 102:19]
    .io_x1(m_91_io_x1),
    .io_x2(m_91_io_x2),
    .io_x3(m_91_io_x3),
    .io_s(m_91_io_s),
    .io_cout(m_91_io_cout)
  );
  Adder m_92 ( // @[MUL.scala 102:19]
    .io_x1(m_92_io_x1),
    .io_x2(m_92_io_x2),
    .io_x3(m_92_io_x3),
    .io_s(m_92_io_s),
    .io_cout(m_92_io_cout)
  );
  Adder m_93 ( // @[MUL.scala 102:19]
    .io_x1(m_93_io_x1),
    .io_x2(m_93_io_x2),
    .io_x3(m_93_io_x3),
    .io_s(m_93_io_s),
    .io_cout(m_93_io_cout)
  );
  Adder m_94 ( // @[MUL.scala 102:19]
    .io_x1(m_94_io_x1),
    .io_x2(m_94_io_x2),
    .io_x3(m_94_io_x3),
    .io_s(m_94_io_s),
    .io_cout(m_94_io_cout)
  );
  Adder m_95 ( // @[MUL.scala 102:19]
    .io_x1(m_95_io_x1),
    .io_x2(m_95_io_x2),
    .io_x3(m_95_io_x3),
    .io_s(m_95_io_s),
    .io_cout(m_95_io_cout)
  );
  Adder m_96 ( // @[MUL.scala 102:19]
    .io_x1(m_96_io_x1),
    .io_x2(m_96_io_x2),
    .io_x3(m_96_io_x3),
    .io_s(m_96_io_s),
    .io_cout(m_96_io_cout)
  );
  Adder m_97 ( // @[MUL.scala 102:19]
    .io_x1(m_97_io_x1),
    .io_x2(m_97_io_x2),
    .io_x3(m_97_io_x3),
    .io_s(m_97_io_s),
    .io_cout(m_97_io_cout)
  );
  Adder m_98 ( // @[MUL.scala 102:19]
    .io_x1(m_98_io_x1),
    .io_x2(m_98_io_x2),
    .io_x3(m_98_io_x3),
    .io_s(m_98_io_s),
    .io_cout(m_98_io_cout)
  );
  Adder m_99 ( // @[MUL.scala 102:19]
    .io_x1(m_99_io_x1),
    .io_x2(m_99_io_x2),
    .io_x3(m_99_io_x3),
    .io_s(m_99_io_s),
    .io_cout(m_99_io_cout)
  );
  Adder m_100 ( // @[MUL.scala 102:19]
    .io_x1(m_100_io_x1),
    .io_x2(m_100_io_x2),
    .io_x3(m_100_io_x3),
    .io_s(m_100_io_s),
    .io_cout(m_100_io_cout)
  );
  Adder m_101 ( // @[MUL.scala 102:19]
    .io_x1(m_101_io_x1),
    .io_x2(m_101_io_x2),
    .io_x3(m_101_io_x3),
    .io_s(m_101_io_s),
    .io_cout(m_101_io_cout)
  );
  Adder m_102 ( // @[MUL.scala 102:19]
    .io_x1(m_102_io_x1),
    .io_x2(m_102_io_x2),
    .io_x3(m_102_io_x3),
    .io_s(m_102_io_s),
    .io_cout(m_102_io_cout)
  );
  Adder m_103 ( // @[MUL.scala 102:19]
    .io_x1(m_103_io_x1),
    .io_x2(m_103_io_x2),
    .io_x3(m_103_io_x3),
    .io_s(m_103_io_s),
    .io_cout(m_103_io_cout)
  );
  Adder m_104 ( // @[MUL.scala 102:19]
    .io_x1(m_104_io_x1),
    .io_x2(m_104_io_x2),
    .io_x3(m_104_io_x3),
    .io_s(m_104_io_s),
    .io_cout(m_104_io_cout)
  );
  Adder m_105 ( // @[MUL.scala 102:19]
    .io_x1(m_105_io_x1),
    .io_x2(m_105_io_x2),
    .io_x3(m_105_io_x3),
    .io_s(m_105_io_s),
    .io_cout(m_105_io_cout)
  );
  Adder m_106 ( // @[MUL.scala 102:19]
    .io_x1(m_106_io_x1),
    .io_x2(m_106_io_x2),
    .io_x3(m_106_io_x3),
    .io_s(m_106_io_s),
    .io_cout(m_106_io_cout)
  );
  Adder m_107 ( // @[MUL.scala 102:19]
    .io_x1(m_107_io_x1),
    .io_x2(m_107_io_x2),
    .io_x3(m_107_io_x3),
    .io_s(m_107_io_s),
    .io_cout(m_107_io_cout)
  );
  Adder m_108 ( // @[MUL.scala 102:19]
    .io_x1(m_108_io_x1),
    .io_x2(m_108_io_x2),
    .io_x3(m_108_io_x3),
    .io_s(m_108_io_s),
    .io_cout(m_108_io_cout)
  );
  Adder m_109 ( // @[MUL.scala 102:19]
    .io_x1(m_109_io_x1),
    .io_x2(m_109_io_x2),
    .io_x3(m_109_io_x3),
    .io_s(m_109_io_s),
    .io_cout(m_109_io_cout)
  );
  Adder m_110 ( // @[MUL.scala 102:19]
    .io_x1(m_110_io_x1),
    .io_x2(m_110_io_x2),
    .io_x3(m_110_io_x3),
    .io_s(m_110_io_s),
    .io_cout(m_110_io_cout)
  );
  Adder m_111 ( // @[MUL.scala 102:19]
    .io_x1(m_111_io_x1),
    .io_x2(m_111_io_x2),
    .io_x3(m_111_io_x3),
    .io_s(m_111_io_s),
    .io_cout(m_111_io_cout)
  );
  Half_Adder m_112 ( // @[MUL.scala 124:19]
    .io_in_0(m_112_io_in_0),
    .io_in_1(m_112_io_in_1),
    .io_out_0(m_112_io_out_0),
    .io_out_1(m_112_io_out_1)
  );
  Adder m_113 ( // @[MUL.scala 102:19]
    .io_x1(m_113_io_x1),
    .io_x2(m_113_io_x2),
    .io_x3(m_113_io_x3),
    .io_s(m_113_io_s),
    .io_cout(m_113_io_cout)
  );
  Adder m_114 ( // @[MUL.scala 102:19]
    .io_x1(m_114_io_x1),
    .io_x2(m_114_io_x2),
    .io_x3(m_114_io_x3),
    .io_s(m_114_io_s),
    .io_cout(m_114_io_cout)
  );
  Adder m_115 ( // @[MUL.scala 102:19]
    .io_x1(m_115_io_x1),
    .io_x2(m_115_io_x2),
    .io_x3(m_115_io_x3),
    .io_s(m_115_io_s),
    .io_cout(m_115_io_cout)
  );
  Adder m_116 ( // @[MUL.scala 102:19]
    .io_x1(m_116_io_x1),
    .io_x2(m_116_io_x2),
    .io_x3(m_116_io_x3),
    .io_s(m_116_io_s),
    .io_cout(m_116_io_cout)
  );
  Adder m_117 ( // @[MUL.scala 102:19]
    .io_x1(m_117_io_x1),
    .io_x2(m_117_io_x2),
    .io_x3(m_117_io_x3),
    .io_s(m_117_io_s),
    .io_cout(m_117_io_cout)
  );
  Half_Adder m_118 ( // @[MUL.scala 124:19]
    .io_in_0(m_118_io_in_0),
    .io_in_1(m_118_io_in_1),
    .io_out_0(m_118_io_out_0),
    .io_out_1(m_118_io_out_1)
  );
  Adder m_119 ( // @[MUL.scala 102:19]
    .io_x1(m_119_io_x1),
    .io_x2(m_119_io_x2),
    .io_x3(m_119_io_x3),
    .io_s(m_119_io_s),
    .io_cout(m_119_io_cout)
  );
  Adder m_120 ( // @[MUL.scala 102:19]
    .io_x1(m_120_io_x1),
    .io_x2(m_120_io_x2),
    .io_x3(m_120_io_x3),
    .io_s(m_120_io_s),
    .io_cout(m_120_io_cout)
  );
  Adder m_121 ( // @[MUL.scala 102:19]
    .io_x1(m_121_io_x1),
    .io_x2(m_121_io_x2),
    .io_x3(m_121_io_x3),
    .io_s(m_121_io_s),
    .io_cout(m_121_io_cout)
  );
  Adder m_122 ( // @[MUL.scala 102:19]
    .io_x1(m_122_io_x1),
    .io_x2(m_122_io_x2),
    .io_x3(m_122_io_x3),
    .io_s(m_122_io_s),
    .io_cout(m_122_io_cout)
  );
  Adder m_123 ( // @[MUL.scala 102:19]
    .io_x1(m_123_io_x1),
    .io_x2(m_123_io_x2),
    .io_x3(m_123_io_x3),
    .io_s(m_123_io_s),
    .io_cout(m_123_io_cout)
  );
  Half_Adder m_124 ( // @[MUL.scala 124:19]
    .io_in_0(m_124_io_in_0),
    .io_in_1(m_124_io_in_1),
    .io_out_0(m_124_io_out_0),
    .io_out_1(m_124_io_out_1)
  );
  Adder m_125 ( // @[MUL.scala 102:19]
    .io_x1(m_125_io_x1),
    .io_x2(m_125_io_x2),
    .io_x3(m_125_io_x3),
    .io_s(m_125_io_s),
    .io_cout(m_125_io_cout)
  );
  Adder m_126 ( // @[MUL.scala 102:19]
    .io_x1(m_126_io_x1),
    .io_x2(m_126_io_x2),
    .io_x3(m_126_io_x3),
    .io_s(m_126_io_s),
    .io_cout(m_126_io_cout)
  );
  Adder m_127 ( // @[MUL.scala 102:19]
    .io_x1(m_127_io_x1),
    .io_x2(m_127_io_x2),
    .io_x3(m_127_io_x3),
    .io_s(m_127_io_s),
    .io_cout(m_127_io_cout)
  );
  Adder m_128 ( // @[MUL.scala 102:19]
    .io_x1(m_128_io_x1),
    .io_x2(m_128_io_x2),
    .io_x3(m_128_io_x3),
    .io_s(m_128_io_s),
    .io_cout(m_128_io_cout)
  );
  Adder m_129 ( // @[MUL.scala 102:19]
    .io_x1(m_129_io_x1),
    .io_x2(m_129_io_x2),
    .io_x3(m_129_io_x3),
    .io_s(m_129_io_s),
    .io_cout(m_129_io_cout)
  );
  Half_Adder m_130 ( // @[MUL.scala 124:19]
    .io_in_0(m_130_io_in_0),
    .io_in_1(m_130_io_in_1),
    .io_out_0(m_130_io_out_0),
    .io_out_1(m_130_io_out_1)
  );
  Adder m_131 ( // @[MUL.scala 102:19]
    .io_x1(m_131_io_x1),
    .io_x2(m_131_io_x2),
    .io_x3(m_131_io_x3),
    .io_s(m_131_io_s),
    .io_cout(m_131_io_cout)
  );
  Adder m_132 ( // @[MUL.scala 102:19]
    .io_x1(m_132_io_x1),
    .io_x2(m_132_io_x2),
    .io_x3(m_132_io_x3),
    .io_s(m_132_io_s),
    .io_cout(m_132_io_cout)
  );
  Adder m_133 ( // @[MUL.scala 102:19]
    .io_x1(m_133_io_x1),
    .io_x2(m_133_io_x2),
    .io_x3(m_133_io_x3),
    .io_s(m_133_io_s),
    .io_cout(m_133_io_cout)
  );
  Adder m_134 ( // @[MUL.scala 102:19]
    .io_x1(m_134_io_x1),
    .io_x2(m_134_io_x2),
    .io_x3(m_134_io_x3),
    .io_s(m_134_io_s),
    .io_cout(m_134_io_cout)
  );
  Adder m_135 ( // @[MUL.scala 102:19]
    .io_x1(m_135_io_x1),
    .io_x2(m_135_io_x2),
    .io_x3(m_135_io_x3),
    .io_s(m_135_io_s),
    .io_cout(m_135_io_cout)
  );
  Half_Adder m_136 ( // @[MUL.scala 124:19]
    .io_in_0(m_136_io_in_0),
    .io_in_1(m_136_io_in_1),
    .io_out_0(m_136_io_out_0),
    .io_out_1(m_136_io_out_1)
  );
  Adder m_137 ( // @[MUL.scala 102:19]
    .io_x1(m_137_io_x1),
    .io_x2(m_137_io_x2),
    .io_x3(m_137_io_x3),
    .io_s(m_137_io_s),
    .io_cout(m_137_io_cout)
  );
  Adder m_138 ( // @[MUL.scala 102:19]
    .io_x1(m_138_io_x1),
    .io_x2(m_138_io_x2),
    .io_x3(m_138_io_x3),
    .io_s(m_138_io_s),
    .io_cout(m_138_io_cout)
  );
  Adder m_139 ( // @[MUL.scala 102:19]
    .io_x1(m_139_io_x1),
    .io_x2(m_139_io_x2),
    .io_x3(m_139_io_x3),
    .io_s(m_139_io_s),
    .io_cout(m_139_io_cout)
  );
  Adder m_140 ( // @[MUL.scala 102:19]
    .io_x1(m_140_io_x1),
    .io_x2(m_140_io_x2),
    .io_x3(m_140_io_x3),
    .io_s(m_140_io_s),
    .io_cout(m_140_io_cout)
  );
  Adder m_141 ( // @[MUL.scala 102:19]
    .io_x1(m_141_io_x1),
    .io_x2(m_141_io_x2),
    .io_x3(m_141_io_x3),
    .io_s(m_141_io_s),
    .io_cout(m_141_io_cout)
  );
  Half_Adder m_142 ( // @[MUL.scala 124:19]
    .io_in_0(m_142_io_in_0),
    .io_in_1(m_142_io_in_1),
    .io_out_0(m_142_io_out_0),
    .io_out_1(m_142_io_out_1)
  );
  Adder m_143 ( // @[MUL.scala 102:19]
    .io_x1(m_143_io_x1),
    .io_x2(m_143_io_x2),
    .io_x3(m_143_io_x3),
    .io_s(m_143_io_s),
    .io_cout(m_143_io_cout)
  );
  Adder m_144 ( // @[MUL.scala 102:19]
    .io_x1(m_144_io_x1),
    .io_x2(m_144_io_x2),
    .io_x3(m_144_io_x3),
    .io_s(m_144_io_s),
    .io_cout(m_144_io_cout)
  );
  Adder m_145 ( // @[MUL.scala 102:19]
    .io_x1(m_145_io_x1),
    .io_x2(m_145_io_x2),
    .io_x3(m_145_io_x3),
    .io_s(m_145_io_s),
    .io_cout(m_145_io_cout)
  );
  Adder m_146 ( // @[MUL.scala 102:19]
    .io_x1(m_146_io_x1),
    .io_x2(m_146_io_x2),
    .io_x3(m_146_io_x3),
    .io_s(m_146_io_s),
    .io_cout(m_146_io_cout)
  );
  Adder m_147 ( // @[MUL.scala 102:19]
    .io_x1(m_147_io_x1),
    .io_x2(m_147_io_x2),
    .io_x3(m_147_io_x3),
    .io_s(m_147_io_s),
    .io_cout(m_147_io_cout)
  );
  Half_Adder m_148 ( // @[MUL.scala 124:19]
    .io_in_0(m_148_io_in_0),
    .io_in_1(m_148_io_in_1),
    .io_out_0(m_148_io_out_0),
    .io_out_1(m_148_io_out_1)
  );
  Adder m_149 ( // @[MUL.scala 102:19]
    .io_x1(m_149_io_x1),
    .io_x2(m_149_io_x2),
    .io_x3(m_149_io_x3),
    .io_s(m_149_io_s),
    .io_cout(m_149_io_cout)
  );
  Adder m_150 ( // @[MUL.scala 102:19]
    .io_x1(m_150_io_x1),
    .io_x2(m_150_io_x2),
    .io_x3(m_150_io_x3),
    .io_s(m_150_io_s),
    .io_cout(m_150_io_cout)
  );
  Adder m_151 ( // @[MUL.scala 102:19]
    .io_x1(m_151_io_x1),
    .io_x2(m_151_io_x2),
    .io_x3(m_151_io_x3),
    .io_s(m_151_io_s),
    .io_cout(m_151_io_cout)
  );
  Adder m_152 ( // @[MUL.scala 102:19]
    .io_x1(m_152_io_x1),
    .io_x2(m_152_io_x2),
    .io_x3(m_152_io_x3),
    .io_s(m_152_io_s),
    .io_cout(m_152_io_cout)
  );
  Adder m_153 ( // @[MUL.scala 102:19]
    .io_x1(m_153_io_x1),
    .io_x2(m_153_io_x2),
    .io_x3(m_153_io_x3),
    .io_s(m_153_io_s),
    .io_cout(m_153_io_cout)
  );
  Adder m_154 ( // @[MUL.scala 102:19]
    .io_x1(m_154_io_x1),
    .io_x2(m_154_io_x2),
    .io_x3(m_154_io_x3),
    .io_s(m_154_io_s),
    .io_cout(m_154_io_cout)
  );
  Adder m_155 ( // @[MUL.scala 102:19]
    .io_x1(m_155_io_x1),
    .io_x2(m_155_io_x2),
    .io_x3(m_155_io_x3),
    .io_s(m_155_io_s),
    .io_cout(m_155_io_cout)
  );
  Adder m_156 ( // @[MUL.scala 102:19]
    .io_x1(m_156_io_x1),
    .io_x2(m_156_io_x2),
    .io_x3(m_156_io_x3),
    .io_s(m_156_io_s),
    .io_cout(m_156_io_cout)
  );
  Adder m_157 ( // @[MUL.scala 102:19]
    .io_x1(m_157_io_x1),
    .io_x2(m_157_io_x2),
    .io_x3(m_157_io_x3),
    .io_s(m_157_io_s),
    .io_cout(m_157_io_cout)
  );
  Adder m_158 ( // @[MUL.scala 102:19]
    .io_x1(m_158_io_x1),
    .io_x2(m_158_io_x2),
    .io_x3(m_158_io_x3),
    .io_s(m_158_io_s),
    .io_cout(m_158_io_cout)
  );
  Adder m_159 ( // @[MUL.scala 102:19]
    .io_x1(m_159_io_x1),
    .io_x2(m_159_io_x2),
    .io_x3(m_159_io_x3),
    .io_s(m_159_io_s),
    .io_cout(m_159_io_cout)
  );
  Adder m_160 ( // @[MUL.scala 102:19]
    .io_x1(m_160_io_x1),
    .io_x2(m_160_io_x2),
    .io_x3(m_160_io_x3),
    .io_s(m_160_io_s),
    .io_cout(m_160_io_cout)
  );
  Adder m_161 ( // @[MUL.scala 102:19]
    .io_x1(m_161_io_x1),
    .io_x2(m_161_io_x2),
    .io_x3(m_161_io_x3),
    .io_s(m_161_io_s),
    .io_cout(m_161_io_cout)
  );
  Adder m_162 ( // @[MUL.scala 102:19]
    .io_x1(m_162_io_x1),
    .io_x2(m_162_io_x2),
    .io_x3(m_162_io_x3),
    .io_s(m_162_io_s),
    .io_cout(m_162_io_cout)
  );
  Adder m_163 ( // @[MUL.scala 102:19]
    .io_x1(m_163_io_x1),
    .io_x2(m_163_io_x2),
    .io_x3(m_163_io_x3),
    .io_s(m_163_io_s),
    .io_cout(m_163_io_cout)
  );
  Adder m_164 ( // @[MUL.scala 102:19]
    .io_x1(m_164_io_x1),
    .io_x2(m_164_io_x2),
    .io_x3(m_164_io_x3),
    .io_s(m_164_io_s),
    .io_cout(m_164_io_cout)
  );
  Adder m_165 ( // @[MUL.scala 102:19]
    .io_x1(m_165_io_x1),
    .io_x2(m_165_io_x2),
    .io_x3(m_165_io_x3),
    .io_s(m_165_io_s),
    .io_cout(m_165_io_cout)
  );
  Adder m_166 ( // @[MUL.scala 102:19]
    .io_x1(m_166_io_x1),
    .io_x2(m_166_io_x2),
    .io_x3(m_166_io_x3),
    .io_s(m_166_io_s),
    .io_cout(m_166_io_cout)
  );
  Adder m_167 ( // @[MUL.scala 102:19]
    .io_x1(m_167_io_x1),
    .io_x2(m_167_io_x2),
    .io_x3(m_167_io_x3),
    .io_s(m_167_io_s),
    .io_cout(m_167_io_cout)
  );
  Half_Adder m_168 ( // @[MUL.scala 124:19]
    .io_in_0(m_168_io_in_0),
    .io_in_1(m_168_io_in_1),
    .io_out_0(m_168_io_out_0),
    .io_out_1(m_168_io_out_1)
  );
  Adder m_169 ( // @[MUL.scala 102:19]
    .io_x1(m_169_io_x1),
    .io_x2(m_169_io_x2),
    .io_x3(m_169_io_x3),
    .io_s(m_169_io_s),
    .io_cout(m_169_io_cout)
  );
  Adder m_170 ( // @[MUL.scala 102:19]
    .io_x1(m_170_io_x1),
    .io_x2(m_170_io_x2),
    .io_x3(m_170_io_x3),
    .io_s(m_170_io_s),
    .io_cout(m_170_io_cout)
  );
  Adder m_171 ( // @[MUL.scala 102:19]
    .io_x1(m_171_io_x1),
    .io_x2(m_171_io_x2),
    .io_x3(m_171_io_x3),
    .io_s(m_171_io_s),
    .io_cout(m_171_io_cout)
  );
  Adder m_172 ( // @[MUL.scala 102:19]
    .io_x1(m_172_io_x1),
    .io_x2(m_172_io_x2),
    .io_x3(m_172_io_x3),
    .io_s(m_172_io_s),
    .io_cout(m_172_io_cout)
  );
  Half_Adder m_173 ( // @[MUL.scala 124:19]
    .io_in_0(m_173_io_in_0),
    .io_in_1(m_173_io_in_1),
    .io_out_0(m_173_io_out_0),
    .io_out_1(m_173_io_out_1)
  );
  Adder m_174 ( // @[MUL.scala 102:19]
    .io_x1(m_174_io_x1),
    .io_x2(m_174_io_x2),
    .io_x3(m_174_io_x3),
    .io_s(m_174_io_s),
    .io_cout(m_174_io_cout)
  );
  Adder m_175 ( // @[MUL.scala 102:19]
    .io_x1(m_175_io_x1),
    .io_x2(m_175_io_x2),
    .io_x3(m_175_io_x3),
    .io_s(m_175_io_s),
    .io_cout(m_175_io_cout)
  );
  Adder m_176 ( // @[MUL.scala 102:19]
    .io_x1(m_176_io_x1),
    .io_x2(m_176_io_x2),
    .io_x3(m_176_io_x3),
    .io_s(m_176_io_s),
    .io_cout(m_176_io_cout)
  );
  Adder m_177 ( // @[MUL.scala 102:19]
    .io_x1(m_177_io_x1),
    .io_x2(m_177_io_x2),
    .io_x3(m_177_io_x3),
    .io_s(m_177_io_s),
    .io_cout(m_177_io_cout)
  );
  Adder m_178 ( // @[MUL.scala 102:19]
    .io_x1(m_178_io_x1),
    .io_x2(m_178_io_x2),
    .io_x3(m_178_io_x3),
    .io_s(m_178_io_s),
    .io_cout(m_178_io_cout)
  );
  Adder m_179 ( // @[MUL.scala 102:19]
    .io_x1(m_179_io_x1),
    .io_x2(m_179_io_x2),
    .io_x3(m_179_io_x3),
    .io_s(m_179_io_s),
    .io_cout(m_179_io_cout)
  );
  Adder m_180 ( // @[MUL.scala 102:19]
    .io_x1(m_180_io_x1),
    .io_x2(m_180_io_x2),
    .io_x3(m_180_io_x3),
    .io_s(m_180_io_s),
    .io_cout(m_180_io_cout)
  );
  Adder m_181 ( // @[MUL.scala 102:19]
    .io_x1(m_181_io_x1),
    .io_x2(m_181_io_x2),
    .io_x3(m_181_io_x3),
    .io_s(m_181_io_s),
    .io_cout(m_181_io_cout)
  );
  Adder m_182 ( // @[MUL.scala 102:19]
    .io_x1(m_182_io_x1),
    .io_x2(m_182_io_x2),
    .io_x3(m_182_io_x3),
    .io_s(m_182_io_s),
    .io_cout(m_182_io_cout)
  );
  Adder m_183 ( // @[MUL.scala 102:19]
    .io_x1(m_183_io_x1),
    .io_x2(m_183_io_x2),
    .io_x3(m_183_io_x3),
    .io_s(m_183_io_s),
    .io_cout(m_183_io_cout)
  );
  Adder m_184 ( // @[MUL.scala 102:19]
    .io_x1(m_184_io_x1),
    .io_x2(m_184_io_x2),
    .io_x3(m_184_io_x3),
    .io_s(m_184_io_s),
    .io_cout(m_184_io_cout)
  );
  Adder m_185 ( // @[MUL.scala 102:19]
    .io_x1(m_185_io_x1),
    .io_x2(m_185_io_x2),
    .io_x3(m_185_io_x3),
    .io_s(m_185_io_s),
    .io_cout(m_185_io_cout)
  );
  Adder m_186 ( // @[MUL.scala 102:19]
    .io_x1(m_186_io_x1),
    .io_x2(m_186_io_x2),
    .io_x3(m_186_io_x3),
    .io_s(m_186_io_s),
    .io_cout(m_186_io_cout)
  );
  Adder m_187 ( // @[MUL.scala 102:19]
    .io_x1(m_187_io_x1),
    .io_x2(m_187_io_x2),
    .io_x3(m_187_io_x3),
    .io_s(m_187_io_s),
    .io_cout(m_187_io_cout)
  );
  Adder m_188 ( // @[MUL.scala 102:19]
    .io_x1(m_188_io_x1),
    .io_x2(m_188_io_x2),
    .io_x3(m_188_io_x3),
    .io_s(m_188_io_s),
    .io_cout(m_188_io_cout)
  );
  Adder m_189 ( // @[MUL.scala 102:19]
    .io_x1(m_189_io_x1),
    .io_x2(m_189_io_x2),
    .io_x3(m_189_io_x3),
    .io_s(m_189_io_s),
    .io_cout(m_189_io_cout)
  );
  Adder m_190 ( // @[MUL.scala 102:19]
    .io_x1(m_190_io_x1),
    .io_x2(m_190_io_x2),
    .io_x3(m_190_io_x3),
    .io_s(m_190_io_s),
    .io_cout(m_190_io_cout)
  );
  Adder m_191 ( // @[MUL.scala 102:19]
    .io_x1(m_191_io_x1),
    .io_x2(m_191_io_x2),
    .io_x3(m_191_io_x3),
    .io_s(m_191_io_s),
    .io_cout(m_191_io_cout)
  );
  Adder m_192 ( // @[MUL.scala 102:19]
    .io_x1(m_192_io_x1),
    .io_x2(m_192_io_x2),
    .io_x3(m_192_io_x3),
    .io_s(m_192_io_s),
    .io_cout(m_192_io_cout)
  );
  Half_Adder m_193 ( // @[MUL.scala 124:19]
    .io_in_0(m_193_io_in_0),
    .io_in_1(m_193_io_in_1),
    .io_out_0(m_193_io_out_0),
    .io_out_1(m_193_io_out_1)
  );
  Adder m_194 ( // @[MUL.scala 102:19]
    .io_x1(m_194_io_x1),
    .io_x2(m_194_io_x2),
    .io_x3(m_194_io_x3),
    .io_s(m_194_io_s),
    .io_cout(m_194_io_cout)
  );
  Adder m_195 ( // @[MUL.scala 102:19]
    .io_x1(m_195_io_x1),
    .io_x2(m_195_io_x2),
    .io_x3(m_195_io_x3),
    .io_s(m_195_io_s),
    .io_cout(m_195_io_cout)
  );
  Adder m_196 ( // @[MUL.scala 102:19]
    .io_x1(m_196_io_x1),
    .io_x2(m_196_io_x2),
    .io_x3(m_196_io_x3),
    .io_s(m_196_io_s),
    .io_cout(m_196_io_cout)
  );
  Half_Adder m_197 ( // @[MUL.scala 124:19]
    .io_in_0(m_197_io_in_0),
    .io_in_1(m_197_io_in_1),
    .io_out_0(m_197_io_out_0),
    .io_out_1(m_197_io_out_1)
  );
  Adder m_198 ( // @[MUL.scala 102:19]
    .io_x1(m_198_io_x1),
    .io_x2(m_198_io_x2),
    .io_x3(m_198_io_x3),
    .io_s(m_198_io_s),
    .io_cout(m_198_io_cout)
  );
  Adder m_199 ( // @[MUL.scala 102:19]
    .io_x1(m_199_io_x1),
    .io_x2(m_199_io_x2),
    .io_x3(m_199_io_x3),
    .io_s(m_199_io_s),
    .io_cout(m_199_io_cout)
  );
  Adder m_200 ( // @[MUL.scala 102:19]
    .io_x1(m_200_io_x1),
    .io_x2(m_200_io_x2),
    .io_x3(m_200_io_x3),
    .io_s(m_200_io_s),
    .io_cout(m_200_io_cout)
  );
  Adder m_201 ( // @[MUL.scala 102:19]
    .io_x1(m_201_io_x1),
    .io_x2(m_201_io_x2),
    .io_x3(m_201_io_x3),
    .io_s(m_201_io_s),
    .io_cout(m_201_io_cout)
  );
  Adder m_202 ( // @[MUL.scala 102:19]
    .io_x1(m_202_io_x1),
    .io_x2(m_202_io_x2),
    .io_x3(m_202_io_x3),
    .io_s(m_202_io_s),
    .io_cout(m_202_io_cout)
  );
  Adder m_203 ( // @[MUL.scala 102:19]
    .io_x1(m_203_io_x1),
    .io_x2(m_203_io_x2),
    .io_x3(m_203_io_x3),
    .io_s(m_203_io_s),
    .io_cout(m_203_io_cout)
  );
  Adder m_204 ( // @[MUL.scala 102:19]
    .io_x1(m_204_io_x1),
    .io_x2(m_204_io_x2),
    .io_x3(m_204_io_x3),
    .io_s(m_204_io_s),
    .io_cout(m_204_io_cout)
  );
  Adder m_205 ( // @[MUL.scala 102:19]
    .io_x1(m_205_io_x1),
    .io_x2(m_205_io_x2),
    .io_x3(m_205_io_x3),
    .io_s(m_205_io_s),
    .io_cout(m_205_io_cout)
  );
  Adder m_206 ( // @[MUL.scala 102:19]
    .io_x1(m_206_io_x1),
    .io_x2(m_206_io_x2),
    .io_x3(m_206_io_x3),
    .io_s(m_206_io_s),
    .io_cout(m_206_io_cout)
  );
  Adder m_207 ( // @[MUL.scala 102:19]
    .io_x1(m_207_io_x1),
    .io_x2(m_207_io_x2),
    .io_x3(m_207_io_x3),
    .io_s(m_207_io_s),
    .io_cout(m_207_io_cout)
  );
  Adder m_208 ( // @[MUL.scala 102:19]
    .io_x1(m_208_io_x1),
    .io_x2(m_208_io_x2),
    .io_x3(m_208_io_x3),
    .io_s(m_208_io_s),
    .io_cout(m_208_io_cout)
  );
  Adder m_209 ( // @[MUL.scala 102:19]
    .io_x1(m_209_io_x1),
    .io_x2(m_209_io_x2),
    .io_x3(m_209_io_x3),
    .io_s(m_209_io_s),
    .io_cout(m_209_io_cout)
  );
  Adder m_210 ( // @[MUL.scala 102:19]
    .io_x1(m_210_io_x1),
    .io_x2(m_210_io_x2),
    .io_x3(m_210_io_x3),
    .io_s(m_210_io_s),
    .io_cout(m_210_io_cout)
  );
  Adder m_211 ( // @[MUL.scala 102:19]
    .io_x1(m_211_io_x1),
    .io_x2(m_211_io_x2),
    .io_x3(m_211_io_x3),
    .io_s(m_211_io_s),
    .io_cout(m_211_io_cout)
  );
  Half_Adder m_212 ( // @[MUL.scala 124:19]
    .io_in_0(m_212_io_in_0),
    .io_in_1(m_212_io_in_1),
    .io_out_0(m_212_io_out_0),
    .io_out_1(m_212_io_out_1)
  );
  Adder m_213 ( // @[MUL.scala 102:19]
    .io_x1(m_213_io_x1),
    .io_x2(m_213_io_x2),
    .io_x3(m_213_io_x3),
    .io_s(m_213_io_s),
    .io_cout(m_213_io_cout)
  );
  Adder m_214 ( // @[MUL.scala 102:19]
    .io_x1(m_214_io_x1),
    .io_x2(m_214_io_x2),
    .io_x3(m_214_io_x3),
    .io_s(m_214_io_s),
    .io_cout(m_214_io_cout)
  );
  Half_Adder m_215 ( // @[MUL.scala 124:19]
    .io_in_0(m_215_io_in_0),
    .io_in_1(m_215_io_in_1),
    .io_out_0(m_215_io_out_0),
    .io_out_1(m_215_io_out_1)
  );
  Adder m_216 ( // @[MUL.scala 102:19]
    .io_x1(m_216_io_x1),
    .io_x2(m_216_io_x2),
    .io_x3(m_216_io_x3),
    .io_s(m_216_io_s),
    .io_cout(m_216_io_cout)
  );
  Adder m_217 ( // @[MUL.scala 102:19]
    .io_x1(m_217_io_x1),
    .io_x2(m_217_io_x2),
    .io_x3(m_217_io_x3),
    .io_s(m_217_io_s),
    .io_cout(m_217_io_cout)
  );
  Adder m_218 ( // @[MUL.scala 102:19]
    .io_x1(m_218_io_x1),
    .io_x2(m_218_io_x2),
    .io_x3(m_218_io_x3),
    .io_s(m_218_io_s),
    .io_cout(m_218_io_cout)
  );
  Adder m_219 ( // @[MUL.scala 102:19]
    .io_x1(m_219_io_x1),
    .io_x2(m_219_io_x2),
    .io_x3(m_219_io_x3),
    .io_s(m_219_io_s),
    .io_cout(m_219_io_cout)
  );
  Adder m_220 ( // @[MUL.scala 102:19]
    .io_x1(m_220_io_x1),
    .io_x2(m_220_io_x2),
    .io_x3(m_220_io_x3),
    .io_s(m_220_io_s),
    .io_cout(m_220_io_cout)
  );
  Adder m_221 ( // @[MUL.scala 102:19]
    .io_x1(m_221_io_x1),
    .io_x2(m_221_io_x2),
    .io_x3(m_221_io_x3),
    .io_s(m_221_io_s),
    .io_cout(m_221_io_cout)
  );
  Adder m_222 ( // @[MUL.scala 102:19]
    .io_x1(m_222_io_x1),
    .io_x2(m_222_io_x2),
    .io_x3(m_222_io_x3),
    .io_s(m_222_io_s),
    .io_cout(m_222_io_cout)
  );
  Adder m_223 ( // @[MUL.scala 102:19]
    .io_x1(m_223_io_x1),
    .io_x2(m_223_io_x2),
    .io_x3(m_223_io_x3),
    .io_s(m_223_io_s),
    .io_cout(m_223_io_cout)
  );
  Adder m_224 ( // @[MUL.scala 102:19]
    .io_x1(m_224_io_x1),
    .io_x2(m_224_io_x2),
    .io_x3(m_224_io_x3),
    .io_s(m_224_io_s),
    .io_cout(m_224_io_cout)
  );
  Half_Adder m_225 ( // @[MUL.scala 124:19]
    .io_in_0(m_225_io_in_0),
    .io_in_1(m_225_io_in_1),
    .io_out_0(m_225_io_out_0),
    .io_out_1(m_225_io_out_1)
  );
  Adder m_226 ( // @[MUL.scala 102:19]
    .io_x1(m_226_io_x1),
    .io_x2(m_226_io_x2),
    .io_x3(m_226_io_x3),
    .io_s(m_226_io_s),
    .io_cout(m_226_io_cout)
  );
  Half_Adder m_227 ( // @[MUL.scala 124:19]
    .io_in_0(m_227_io_in_0),
    .io_in_1(m_227_io_in_1),
    .io_out_0(m_227_io_out_0),
    .io_out_1(m_227_io_out_1)
  );
  Adder m_228 ( // @[MUL.scala 102:19]
    .io_x1(m_228_io_x1),
    .io_x2(m_228_io_x2),
    .io_x3(m_228_io_x3),
    .io_s(m_228_io_s),
    .io_cout(m_228_io_cout)
  );
  Adder m_229 ( // @[MUL.scala 102:19]
    .io_x1(m_229_io_x1),
    .io_x2(m_229_io_x2),
    .io_x3(m_229_io_x3),
    .io_s(m_229_io_s),
    .io_cout(m_229_io_cout)
  );
  Adder m_230 ( // @[MUL.scala 102:19]
    .io_x1(m_230_io_x1),
    .io_x2(m_230_io_x2),
    .io_x3(m_230_io_x3),
    .io_s(m_230_io_s),
    .io_cout(m_230_io_cout)
  );
  Adder m_231 ( // @[MUL.scala 102:19]
    .io_x1(m_231_io_x1),
    .io_x2(m_231_io_x2),
    .io_x3(m_231_io_x3),
    .io_s(m_231_io_s),
    .io_cout(m_231_io_cout)
  );
  Half_Adder m_232 ( // @[MUL.scala 124:19]
    .io_in_0(m_232_io_in_0),
    .io_in_1(m_232_io_in_1),
    .io_out_0(m_232_io_out_0),
    .io_out_1(m_232_io_out_1)
  );
  Half_Adder m_233 ( // @[MUL.scala 124:19]
    .io_in_0(m_233_io_in_0),
    .io_in_1(m_233_io_in_1),
    .io_out_0(m_233_io_out_0),
    .io_out_1(m_233_io_out_1)
  );
  Half_Adder m_234 ( // @[MUL.scala 124:19]
    .io_in_0(m_234_io_in_0),
    .io_in_1(m_234_io_in_1),
    .io_out_0(m_234_io_out_0),
    .io_out_1(m_234_io_out_1)
  );
  Half_Adder m_235 ( // @[MUL.scala 124:19]
    .io_in_0(m_235_io_in_0),
    .io_in_1(m_235_io_in_1),
    .io_out_0(m_235_io_out_0),
    .io_out_1(m_235_io_out_1)
  );
  Half_Adder m_236 ( // @[MUL.scala 124:19]
    .io_in_0(m_236_io_in_0),
    .io_in_1(m_236_io_in_1),
    .io_out_0(m_236_io_out_0),
    .io_out_1(m_236_io_out_1)
  );
  Adder m_237 ( // @[MUL.scala 102:19]
    .io_x1(m_237_io_x1),
    .io_x2(m_237_io_x2),
    .io_x3(m_237_io_x3),
    .io_s(m_237_io_s),
    .io_cout(m_237_io_cout)
  );
  Adder m_238 ( // @[MUL.scala 102:19]
    .io_x1(m_238_io_x1),
    .io_x2(m_238_io_x2),
    .io_x3(m_238_io_x3),
    .io_s(m_238_io_s),
    .io_cout(m_238_io_cout)
  );
  Adder m_239 ( // @[MUL.scala 102:19]
    .io_x1(m_239_io_x1),
    .io_x2(m_239_io_x2),
    .io_x3(m_239_io_x3),
    .io_s(m_239_io_s),
    .io_cout(m_239_io_cout)
  );
  Adder m_240 ( // @[MUL.scala 102:19]
    .io_x1(m_240_io_x1),
    .io_x2(m_240_io_x2),
    .io_x3(m_240_io_x3),
    .io_s(m_240_io_s),
    .io_cout(m_240_io_cout)
  );
  Adder m_241 ( // @[MUL.scala 102:19]
    .io_x1(m_241_io_x1),
    .io_x2(m_241_io_x2),
    .io_x3(m_241_io_x3),
    .io_s(m_241_io_s),
    .io_cout(m_241_io_cout)
  );
  Adder m_242 ( // @[MUL.scala 102:19]
    .io_x1(m_242_io_x1),
    .io_x2(m_242_io_x2),
    .io_x3(m_242_io_x3),
    .io_s(m_242_io_s),
    .io_cout(m_242_io_cout)
  );
  Adder m_243 ( // @[MUL.scala 102:19]
    .io_x1(m_243_io_x1),
    .io_x2(m_243_io_x2),
    .io_x3(m_243_io_x3),
    .io_s(m_243_io_s),
    .io_cout(m_243_io_cout)
  );
  Half_Adder m_244 ( // @[MUL.scala 124:19]
    .io_in_0(m_244_io_in_0),
    .io_in_1(m_244_io_in_1),
    .io_out_0(m_244_io_out_0),
    .io_out_1(m_244_io_out_1)
  );
  Adder m_245 ( // @[MUL.scala 102:19]
    .io_x1(m_245_io_x1),
    .io_x2(m_245_io_x2),
    .io_x3(m_245_io_x3),
    .io_s(m_245_io_s),
    .io_cout(m_245_io_cout)
  );
  Half_Adder m_246 ( // @[MUL.scala 124:19]
    .io_in_0(m_246_io_in_0),
    .io_in_1(m_246_io_in_1),
    .io_out_0(m_246_io_out_0),
    .io_out_1(m_246_io_out_1)
  );
  Adder m_247 ( // @[MUL.scala 102:19]
    .io_x1(m_247_io_x1),
    .io_x2(m_247_io_x2),
    .io_x3(m_247_io_x3),
    .io_s(m_247_io_s),
    .io_cout(m_247_io_cout)
  );
  Half_Adder m_248 ( // @[MUL.scala 124:19]
    .io_in_0(m_248_io_in_0),
    .io_in_1(m_248_io_in_1),
    .io_out_0(m_248_io_out_0),
    .io_out_1(m_248_io_out_1)
  );
  Adder m_249 ( // @[MUL.scala 102:19]
    .io_x1(m_249_io_x1),
    .io_x2(m_249_io_x2),
    .io_x3(m_249_io_x3),
    .io_s(m_249_io_s),
    .io_cout(m_249_io_cout)
  );
  Adder m_250 ( // @[MUL.scala 102:19]
    .io_x1(m_250_io_x1),
    .io_x2(m_250_io_x2),
    .io_x3(m_250_io_x3),
    .io_s(m_250_io_s),
    .io_cout(m_250_io_cout)
  );
  Adder m_251 ( // @[MUL.scala 102:19]
    .io_x1(m_251_io_x1),
    .io_x2(m_251_io_x2),
    .io_x3(m_251_io_x3),
    .io_s(m_251_io_s),
    .io_cout(m_251_io_cout)
  );
  Adder m_252 ( // @[MUL.scala 102:19]
    .io_x1(m_252_io_x1),
    .io_x2(m_252_io_x2),
    .io_x3(m_252_io_x3),
    .io_s(m_252_io_s),
    .io_cout(m_252_io_cout)
  );
  Adder m_253 ( // @[MUL.scala 102:19]
    .io_x1(m_253_io_x1),
    .io_x2(m_253_io_x2),
    .io_x3(m_253_io_x3),
    .io_s(m_253_io_s),
    .io_cout(m_253_io_cout)
  );
  Adder m_254 ( // @[MUL.scala 102:19]
    .io_x1(m_254_io_x1),
    .io_x2(m_254_io_x2),
    .io_x3(m_254_io_x3),
    .io_s(m_254_io_s),
    .io_cout(m_254_io_cout)
  );
  Adder m_255 ( // @[MUL.scala 102:19]
    .io_x1(m_255_io_x1),
    .io_x2(m_255_io_x2),
    .io_x3(m_255_io_x3),
    .io_s(m_255_io_s),
    .io_cout(m_255_io_cout)
  );
  Adder m_256 ( // @[MUL.scala 102:19]
    .io_x1(m_256_io_x1),
    .io_x2(m_256_io_x2),
    .io_x3(m_256_io_x3),
    .io_s(m_256_io_s),
    .io_cout(m_256_io_cout)
  );
  Adder m_257 ( // @[MUL.scala 102:19]
    .io_x1(m_257_io_x1),
    .io_x2(m_257_io_x2),
    .io_x3(m_257_io_x3),
    .io_s(m_257_io_s),
    .io_cout(m_257_io_cout)
  );
  Adder m_258 ( // @[MUL.scala 102:19]
    .io_x1(m_258_io_x1),
    .io_x2(m_258_io_x2),
    .io_x3(m_258_io_x3),
    .io_s(m_258_io_s),
    .io_cout(m_258_io_cout)
  );
  Adder m_259 ( // @[MUL.scala 102:19]
    .io_x1(m_259_io_x1),
    .io_x2(m_259_io_x2),
    .io_x3(m_259_io_x3),
    .io_s(m_259_io_s),
    .io_cout(m_259_io_cout)
  );
  Adder m_260 ( // @[MUL.scala 102:19]
    .io_x1(m_260_io_x1),
    .io_x2(m_260_io_x2),
    .io_x3(m_260_io_x3),
    .io_s(m_260_io_s),
    .io_cout(m_260_io_cout)
  );
  Adder m_261 ( // @[MUL.scala 102:19]
    .io_x1(m_261_io_x1),
    .io_x2(m_261_io_x2),
    .io_x3(m_261_io_x3),
    .io_s(m_261_io_s),
    .io_cout(m_261_io_cout)
  );
  Adder m_262 ( // @[MUL.scala 102:19]
    .io_x1(m_262_io_x1),
    .io_x2(m_262_io_x2),
    .io_x3(m_262_io_x3),
    .io_s(m_262_io_s),
    .io_cout(m_262_io_cout)
  );
  Half_Adder m_263 ( // @[MUL.scala 124:19]
    .io_in_0(m_263_io_in_0),
    .io_in_1(m_263_io_in_1),
    .io_out_0(m_263_io_out_0),
    .io_out_1(m_263_io_out_1)
  );
  Adder m_264 ( // @[MUL.scala 102:19]
    .io_x1(m_264_io_x1),
    .io_x2(m_264_io_x2),
    .io_x3(m_264_io_x3),
    .io_s(m_264_io_s),
    .io_cout(m_264_io_cout)
  );
  Adder m_265 ( // @[MUL.scala 102:19]
    .io_x1(m_265_io_x1),
    .io_x2(m_265_io_x2),
    .io_x3(m_265_io_x3),
    .io_s(m_265_io_s),
    .io_cout(m_265_io_cout)
  );
  Half_Adder m_266 ( // @[MUL.scala 124:19]
    .io_in_0(m_266_io_in_0),
    .io_in_1(m_266_io_in_1),
    .io_out_0(m_266_io_out_0),
    .io_out_1(m_266_io_out_1)
  );
  Adder m_267 ( // @[MUL.scala 102:19]
    .io_x1(m_267_io_x1),
    .io_x2(m_267_io_x2),
    .io_x3(m_267_io_x3),
    .io_s(m_267_io_s),
    .io_cout(m_267_io_cout)
  );
  Adder m_268 ( // @[MUL.scala 102:19]
    .io_x1(m_268_io_x1),
    .io_x2(m_268_io_x2),
    .io_x3(m_268_io_x3),
    .io_s(m_268_io_s),
    .io_cout(m_268_io_cout)
  );
  Half_Adder m_269 ( // @[MUL.scala 124:19]
    .io_in_0(m_269_io_in_0),
    .io_in_1(m_269_io_in_1),
    .io_out_0(m_269_io_out_0),
    .io_out_1(m_269_io_out_1)
  );
  Adder m_270 ( // @[MUL.scala 102:19]
    .io_x1(m_270_io_x1),
    .io_x2(m_270_io_x2),
    .io_x3(m_270_io_x3),
    .io_s(m_270_io_s),
    .io_cout(m_270_io_cout)
  );
  Adder m_271 ( // @[MUL.scala 102:19]
    .io_x1(m_271_io_x1),
    .io_x2(m_271_io_x2),
    .io_x3(m_271_io_x3),
    .io_s(m_271_io_s),
    .io_cout(m_271_io_cout)
  );
  Adder m_272 ( // @[MUL.scala 102:19]
    .io_x1(m_272_io_x1),
    .io_x2(m_272_io_x2),
    .io_x3(m_272_io_x3),
    .io_s(m_272_io_s),
    .io_cout(m_272_io_cout)
  );
  Adder m_273 ( // @[MUL.scala 102:19]
    .io_x1(m_273_io_x1),
    .io_x2(m_273_io_x2),
    .io_x3(m_273_io_x3),
    .io_s(m_273_io_s),
    .io_cout(m_273_io_cout)
  );
  Adder m_274 ( // @[MUL.scala 102:19]
    .io_x1(m_274_io_x1),
    .io_x2(m_274_io_x2),
    .io_x3(m_274_io_x3),
    .io_s(m_274_io_s),
    .io_cout(m_274_io_cout)
  );
  Adder m_275 ( // @[MUL.scala 102:19]
    .io_x1(m_275_io_x1),
    .io_x2(m_275_io_x2),
    .io_x3(m_275_io_x3),
    .io_s(m_275_io_s),
    .io_cout(m_275_io_cout)
  );
  Adder m_276 ( // @[MUL.scala 102:19]
    .io_x1(m_276_io_x1),
    .io_x2(m_276_io_x2),
    .io_x3(m_276_io_x3),
    .io_s(m_276_io_s),
    .io_cout(m_276_io_cout)
  );
  Adder m_277 ( // @[MUL.scala 102:19]
    .io_x1(m_277_io_x1),
    .io_x2(m_277_io_x2),
    .io_x3(m_277_io_x3),
    .io_s(m_277_io_s),
    .io_cout(m_277_io_cout)
  );
  Adder m_278 ( // @[MUL.scala 102:19]
    .io_x1(m_278_io_x1),
    .io_x2(m_278_io_x2),
    .io_x3(m_278_io_x3),
    .io_s(m_278_io_s),
    .io_cout(m_278_io_cout)
  );
  Adder m_279 ( // @[MUL.scala 102:19]
    .io_x1(m_279_io_x1),
    .io_x2(m_279_io_x2),
    .io_x3(m_279_io_x3),
    .io_s(m_279_io_s),
    .io_cout(m_279_io_cout)
  );
  Adder m_280 ( // @[MUL.scala 102:19]
    .io_x1(m_280_io_x1),
    .io_x2(m_280_io_x2),
    .io_x3(m_280_io_x3),
    .io_s(m_280_io_s),
    .io_cout(m_280_io_cout)
  );
  Adder m_281 ( // @[MUL.scala 102:19]
    .io_x1(m_281_io_x1),
    .io_x2(m_281_io_x2),
    .io_x3(m_281_io_x3),
    .io_s(m_281_io_s),
    .io_cout(m_281_io_cout)
  );
  Adder m_282 ( // @[MUL.scala 102:19]
    .io_x1(m_282_io_x1),
    .io_x2(m_282_io_x2),
    .io_x3(m_282_io_x3),
    .io_s(m_282_io_s),
    .io_cout(m_282_io_cout)
  );
  Adder m_283 ( // @[MUL.scala 102:19]
    .io_x1(m_283_io_x1),
    .io_x2(m_283_io_x2),
    .io_x3(m_283_io_x3),
    .io_s(m_283_io_s),
    .io_cout(m_283_io_cout)
  );
  Adder m_284 ( // @[MUL.scala 102:19]
    .io_x1(m_284_io_x1),
    .io_x2(m_284_io_x2),
    .io_x3(m_284_io_x3),
    .io_s(m_284_io_s),
    .io_cout(m_284_io_cout)
  );
  Adder m_285 ( // @[MUL.scala 102:19]
    .io_x1(m_285_io_x1),
    .io_x2(m_285_io_x2),
    .io_x3(m_285_io_x3),
    .io_s(m_285_io_s),
    .io_cout(m_285_io_cout)
  );
  Adder m_286 ( // @[MUL.scala 102:19]
    .io_x1(m_286_io_x1),
    .io_x2(m_286_io_x2),
    .io_x3(m_286_io_x3),
    .io_s(m_286_io_s),
    .io_cout(m_286_io_cout)
  );
  Adder m_287 ( // @[MUL.scala 102:19]
    .io_x1(m_287_io_x1),
    .io_x2(m_287_io_x2),
    .io_x3(m_287_io_x3),
    .io_s(m_287_io_s),
    .io_cout(m_287_io_cout)
  );
  Adder m_288 ( // @[MUL.scala 102:19]
    .io_x1(m_288_io_x1),
    .io_x2(m_288_io_x2),
    .io_x3(m_288_io_x3),
    .io_s(m_288_io_s),
    .io_cout(m_288_io_cout)
  );
  Adder m_289 ( // @[MUL.scala 102:19]
    .io_x1(m_289_io_x1),
    .io_x2(m_289_io_x2),
    .io_x3(m_289_io_x3),
    .io_s(m_289_io_s),
    .io_cout(m_289_io_cout)
  );
  Adder m_290 ( // @[MUL.scala 102:19]
    .io_x1(m_290_io_x1),
    .io_x2(m_290_io_x2),
    .io_x3(m_290_io_x3),
    .io_s(m_290_io_s),
    .io_cout(m_290_io_cout)
  );
  Half_Adder m_291 ( // @[MUL.scala 124:19]
    .io_in_0(m_291_io_in_0),
    .io_in_1(m_291_io_in_1),
    .io_out_0(m_291_io_out_0),
    .io_out_1(m_291_io_out_1)
  );
  Adder m_292 ( // @[MUL.scala 102:19]
    .io_x1(m_292_io_x1),
    .io_x2(m_292_io_x2),
    .io_x3(m_292_io_x3),
    .io_s(m_292_io_s),
    .io_cout(m_292_io_cout)
  );
  Adder m_293 ( // @[MUL.scala 102:19]
    .io_x1(m_293_io_x1),
    .io_x2(m_293_io_x2),
    .io_x3(m_293_io_x3),
    .io_s(m_293_io_s),
    .io_cout(m_293_io_cout)
  );
  Adder m_294 ( // @[MUL.scala 102:19]
    .io_x1(m_294_io_x1),
    .io_x2(m_294_io_x2),
    .io_x3(m_294_io_x3),
    .io_s(m_294_io_s),
    .io_cout(m_294_io_cout)
  );
  Half_Adder m_295 ( // @[MUL.scala 124:19]
    .io_in_0(m_295_io_in_0),
    .io_in_1(m_295_io_in_1),
    .io_out_0(m_295_io_out_0),
    .io_out_1(m_295_io_out_1)
  );
  Adder m_296 ( // @[MUL.scala 102:19]
    .io_x1(m_296_io_x1),
    .io_x2(m_296_io_x2),
    .io_x3(m_296_io_x3),
    .io_s(m_296_io_s),
    .io_cout(m_296_io_cout)
  );
  Adder m_297 ( // @[MUL.scala 102:19]
    .io_x1(m_297_io_x1),
    .io_x2(m_297_io_x2),
    .io_x3(m_297_io_x3),
    .io_s(m_297_io_s),
    .io_cout(m_297_io_cout)
  );
  Adder m_298 ( // @[MUL.scala 102:19]
    .io_x1(m_298_io_x1),
    .io_x2(m_298_io_x2),
    .io_x3(m_298_io_x3),
    .io_s(m_298_io_s),
    .io_cout(m_298_io_cout)
  );
  Half_Adder m_299 ( // @[MUL.scala 124:19]
    .io_in_0(m_299_io_in_0),
    .io_in_1(m_299_io_in_1),
    .io_out_0(m_299_io_out_0),
    .io_out_1(m_299_io_out_1)
  );
  Adder m_300 ( // @[MUL.scala 102:19]
    .io_x1(m_300_io_x1),
    .io_x2(m_300_io_x2),
    .io_x3(m_300_io_x3),
    .io_s(m_300_io_s),
    .io_cout(m_300_io_cout)
  );
  Adder m_301 ( // @[MUL.scala 102:19]
    .io_x1(m_301_io_x1),
    .io_x2(m_301_io_x2),
    .io_x3(m_301_io_x3),
    .io_s(m_301_io_s),
    .io_cout(m_301_io_cout)
  );
  Adder m_302 ( // @[MUL.scala 102:19]
    .io_x1(m_302_io_x1),
    .io_x2(m_302_io_x2),
    .io_x3(m_302_io_x3),
    .io_s(m_302_io_s),
    .io_cout(m_302_io_cout)
  );
  Adder m_303 ( // @[MUL.scala 102:19]
    .io_x1(m_303_io_x1),
    .io_x2(m_303_io_x2),
    .io_x3(m_303_io_x3),
    .io_s(m_303_io_s),
    .io_cout(m_303_io_cout)
  );
  Adder m_304 ( // @[MUL.scala 102:19]
    .io_x1(m_304_io_x1),
    .io_x2(m_304_io_x2),
    .io_x3(m_304_io_x3),
    .io_s(m_304_io_s),
    .io_cout(m_304_io_cout)
  );
  Adder m_305 ( // @[MUL.scala 102:19]
    .io_x1(m_305_io_x1),
    .io_x2(m_305_io_x2),
    .io_x3(m_305_io_x3),
    .io_s(m_305_io_s),
    .io_cout(m_305_io_cout)
  );
  Adder m_306 ( // @[MUL.scala 102:19]
    .io_x1(m_306_io_x1),
    .io_x2(m_306_io_x2),
    .io_x3(m_306_io_x3),
    .io_s(m_306_io_s),
    .io_cout(m_306_io_cout)
  );
  Adder m_307 ( // @[MUL.scala 102:19]
    .io_x1(m_307_io_x1),
    .io_x2(m_307_io_x2),
    .io_x3(m_307_io_x3),
    .io_s(m_307_io_s),
    .io_cout(m_307_io_cout)
  );
  Adder m_308 ( // @[MUL.scala 102:19]
    .io_x1(m_308_io_x1),
    .io_x2(m_308_io_x2),
    .io_x3(m_308_io_x3),
    .io_s(m_308_io_s),
    .io_cout(m_308_io_cout)
  );
  Adder m_309 ( // @[MUL.scala 102:19]
    .io_x1(m_309_io_x1),
    .io_x2(m_309_io_x2),
    .io_x3(m_309_io_x3),
    .io_s(m_309_io_s),
    .io_cout(m_309_io_cout)
  );
  Adder m_310 ( // @[MUL.scala 102:19]
    .io_x1(m_310_io_x1),
    .io_x2(m_310_io_x2),
    .io_x3(m_310_io_x3),
    .io_s(m_310_io_s),
    .io_cout(m_310_io_cout)
  );
  Adder m_311 ( // @[MUL.scala 102:19]
    .io_x1(m_311_io_x1),
    .io_x2(m_311_io_x2),
    .io_x3(m_311_io_x3),
    .io_s(m_311_io_s),
    .io_cout(m_311_io_cout)
  );
  Adder m_312 ( // @[MUL.scala 102:19]
    .io_x1(m_312_io_x1),
    .io_x2(m_312_io_x2),
    .io_x3(m_312_io_x3),
    .io_s(m_312_io_s),
    .io_cout(m_312_io_cout)
  );
  Adder m_313 ( // @[MUL.scala 102:19]
    .io_x1(m_313_io_x1),
    .io_x2(m_313_io_x2),
    .io_x3(m_313_io_x3),
    .io_s(m_313_io_s),
    .io_cout(m_313_io_cout)
  );
  Adder m_314 ( // @[MUL.scala 102:19]
    .io_x1(m_314_io_x1),
    .io_x2(m_314_io_x2),
    .io_x3(m_314_io_x3),
    .io_s(m_314_io_s),
    .io_cout(m_314_io_cout)
  );
  Adder m_315 ( // @[MUL.scala 102:19]
    .io_x1(m_315_io_x1),
    .io_x2(m_315_io_x2),
    .io_x3(m_315_io_x3),
    .io_s(m_315_io_s),
    .io_cout(m_315_io_cout)
  );
  Adder m_316 ( // @[MUL.scala 102:19]
    .io_x1(m_316_io_x1),
    .io_x2(m_316_io_x2),
    .io_x3(m_316_io_x3),
    .io_s(m_316_io_s),
    .io_cout(m_316_io_cout)
  );
  Adder m_317 ( // @[MUL.scala 102:19]
    .io_x1(m_317_io_x1),
    .io_x2(m_317_io_x2),
    .io_x3(m_317_io_x3),
    .io_s(m_317_io_s),
    .io_cout(m_317_io_cout)
  );
  Adder m_318 ( // @[MUL.scala 102:19]
    .io_x1(m_318_io_x1),
    .io_x2(m_318_io_x2),
    .io_x3(m_318_io_x3),
    .io_s(m_318_io_s),
    .io_cout(m_318_io_cout)
  );
  Adder m_319 ( // @[MUL.scala 102:19]
    .io_x1(m_319_io_x1),
    .io_x2(m_319_io_x2),
    .io_x3(m_319_io_x3),
    .io_s(m_319_io_s),
    .io_cout(m_319_io_cout)
  );
  Adder m_320 ( // @[MUL.scala 102:19]
    .io_x1(m_320_io_x1),
    .io_x2(m_320_io_x2),
    .io_x3(m_320_io_x3),
    .io_s(m_320_io_s),
    .io_cout(m_320_io_cout)
  );
  Adder m_321 ( // @[MUL.scala 102:19]
    .io_x1(m_321_io_x1),
    .io_x2(m_321_io_x2),
    .io_x3(m_321_io_x3),
    .io_s(m_321_io_s),
    .io_cout(m_321_io_cout)
  );
  Adder m_322 ( // @[MUL.scala 102:19]
    .io_x1(m_322_io_x1),
    .io_x2(m_322_io_x2),
    .io_x3(m_322_io_x3),
    .io_s(m_322_io_s),
    .io_cout(m_322_io_cout)
  );
  Adder m_323 ( // @[MUL.scala 102:19]
    .io_x1(m_323_io_x1),
    .io_x2(m_323_io_x2),
    .io_x3(m_323_io_x3),
    .io_s(m_323_io_s),
    .io_cout(m_323_io_cout)
  );
  Adder m_324 ( // @[MUL.scala 102:19]
    .io_x1(m_324_io_x1),
    .io_x2(m_324_io_x2),
    .io_x3(m_324_io_x3),
    .io_s(m_324_io_s),
    .io_cout(m_324_io_cout)
  );
  Adder m_325 ( // @[MUL.scala 102:19]
    .io_x1(m_325_io_x1),
    .io_x2(m_325_io_x2),
    .io_x3(m_325_io_x3),
    .io_s(m_325_io_s),
    .io_cout(m_325_io_cout)
  );
  Adder m_326 ( // @[MUL.scala 102:19]
    .io_x1(m_326_io_x1),
    .io_x2(m_326_io_x2),
    .io_x3(m_326_io_x3),
    .io_s(m_326_io_s),
    .io_cout(m_326_io_cout)
  );
  Adder m_327 ( // @[MUL.scala 102:19]
    .io_x1(m_327_io_x1),
    .io_x2(m_327_io_x2),
    .io_x3(m_327_io_x3),
    .io_s(m_327_io_s),
    .io_cout(m_327_io_cout)
  );
  Adder m_328 ( // @[MUL.scala 102:19]
    .io_x1(m_328_io_x1),
    .io_x2(m_328_io_x2),
    .io_x3(m_328_io_x3),
    .io_s(m_328_io_s),
    .io_cout(m_328_io_cout)
  );
  Adder m_329 ( // @[MUL.scala 102:19]
    .io_x1(m_329_io_x1),
    .io_x2(m_329_io_x2),
    .io_x3(m_329_io_x3),
    .io_s(m_329_io_s),
    .io_cout(m_329_io_cout)
  );
  Adder m_330 ( // @[MUL.scala 102:19]
    .io_x1(m_330_io_x1),
    .io_x2(m_330_io_x2),
    .io_x3(m_330_io_x3),
    .io_s(m_330_io_s),
    .io_cout(m_330_io_cout)
  );
  Adder m_331 ( // @[MUL.scala 102:19]
    .io_x1(m_331_io_x1),
    .io_x2(m_331_io_x2),
    .io_x3(m_331_io_x3),
    .io_s(m_331_io_s),
    .io_cout(m_331_io_cout)
  );
  Adder m_332 ( // @[MUL.scala 102:19]
    .io_x1(m_332_io_x1),
    .io_x2(m_332_io_x2),
    .io_x3(m_332_io_x3),
    .io_s(m_332_io_s),
    .io_cout(m_332_io_cout)
  );
  Adder m_333 ( // @[MUL.scala 102:19]
    .io_x1(m_333_io_x1),
    .io_x2(m_333_io_x2),
    .io_x3(m_333_io_x3),
    .io_s(m_333_io_s),
    .io_cout(m_333_io_cout)
  );
  Adder m_334 ( // @[MUL.scala 102:19]
    .io_x1(m_334_io_x1),
    .io_x2(m_334_io_x2),
    .io_x3(m_334_io_x3),
    .io_s(m_334_io_s),
    .io_cout(m_334_io_cout)
  );
  Adder m_335 ( // @[MUL.scala 102:19]
    .io_x1(m_335_io_x1),
    .io_x2(m_335_io_x2),
    .io_x3(m_335_io_x3),
    .io_s(m_335_io_s),
    .io_cout(m_335_io_cout)
  );
  Adder m_336 ( // @[MUL.scala 102:19]
    .io_x1(m_336_io_x1),
    .io_x2(m_336_io_x2),
    .io_x3(m_336_io_x3),
    .io_s(m_336_io_s),
    .io_cout(m_336_io_cout)
  );
  Adder m_337 ( // @[MUL.scala 102:19]
    .io_x1(m_337_io_x1),
    .io_x2(m_337_io_x2),
    .io_x3(m_337_io_x3),
    .io_s(m_337_io_s),
    .io_cout(m_337_io_cout)
  );
  Adder m_338 ( // @[MUL.scala 102:19]
    .io_x1(m_338_io_x1),
    .io_x2(m_338_io_x2),
    .io_x3(m_338_io_x3),
    .io_s(m_338_io_s),
    .io_cout(m_338_io_cout)
  );
  Adder m_339 ( // @[MUL.scala 102:19]
    .io_x1(m_339_io_x1),
    .io_x2(m_339_io_x2),
    .io_x3(m_339_io_x3),
    .io_s(m_339_io_s),
    .io_cout(m_339_io_cout)
  );
  Adder m_340 ( // @[MUL.scala 102:19]
    .io_x1(m_340_io_x1),
    .io_x2(m_340_io_x2),
    .io_x3(m_340_io_x3),
    .io_s(m_340_io_s),
    .io_cout(m_340_io_cout)
  );
  Adder m_341 ( // @[MUL.scala 102:19]
    .io_x1(m_341_io_x1),
    .io_x2(m_341_io_x2),
    .io_x3(m_341_io_x3),
    .io_s(m_341_io_s),
    .io_cout(m_341_io_cout)
  );
  Adder m_342 ( // @[MUL.scala 102:19]
    .io_x1(m_342_io_x1),
    .io_x2(m_342_io_x2),
    .io_x3(m_342_io_x3),
    .io_s(m_342_io_s),
    .io_cout(m_342_io_cout)
  );
  Adder m_343 ( // @[MUL.scala 102:19]
    .io_x1(m_343_io_x1),
    .io_x2(m_343_io_x2),
    .io_x3(m_343_io_x3),
    .io_s(m_343_io_s),
    .io_cout(m_343_io_cout)
  );
  Adder m_344 ( // @[MUL.scala 102:19]
    .io_x1(m_344_io_x1),
    .io_x2(m_344_io_x2),
    .io_x3(m_344_io_x3),
    .io_s(m_344_io_s),
    .io_cout(m_344_io_cout)
  );
  Adder m_345 ( // @[MUL.scala 102:19]
    .io_x1(m_345_io_x1),
    .io_x2(m_345_io_x2),
    .io_x3(m_345_io_x3),
    .io_s(m_345_io_s),
    .io_cout(m_345_io_cout)
  );
  Adder m_346 ( // @[MUL.scala 102:19]
    .io_x1(m_346_io_x1),
    .io_x2(m_346_io_x2),
    .io_x3(m_346_io_x3),
    .io_s(m_346_io_s),
    .io_cout(m_346_io_cout)
  );
  Adder m_347 ( // @[MUL.scala 102:19]
    .io_x1(m_347_io_x1),
    .io_x2(m_347_io_x2),
    .io_x3(m_347_io_x3),
    .io_s(m_347_io_s),
    .io_cout(m_347_io_cout)
  );
  Half_Adder m_348 ( // @[MUL.scala 124:19]
    .io_in_0(m_348_io_in_0),
    .io_in_1(m_348_io_in_1),
    .io_out_0(m_348_io_out_0),
    .io_out_1(m_348_io_out_1)
  );
  Adder m_349 ( // @[MUL.scala 102:19]
    .io_x1(m_349_io_x1),
    .io_x2(m_349_io_x2),
    .io_x3(m_349_io_x3),
    .io_s(m_349_io_s),
    .io_cout(m_349_io_cout)
  );
  Adder m_350 ( // @[MUL.scala 102:19]
    .io_x1(m_350_io_x1),
    .io_x2(m_350_io_x2),
    .io_x3(m_350_io_x3),
    .io_s(m_350_io_s),
    .io_cout(m_350_io_cout)
  );
  Half_Adder m_351 ( // @[MUL.scala 124:19]
    .io_in_0(m_351_io_in_0),
    .io_in_1(m_351_io_in_1),
    .io_out_0(m_351_io_out_0),
    .io_out_1(m_351_io_out_1)
  );
  Adder m_352 ( // @[MUL.scala 102:19]
    .io_x1(m_352_io_x1),
    .io_x2(m_352_io_x2),
    .io_x3(m_352_io_x3),
    .io_s(m_352_io_s),
    .io_cout(m_352_io_cout)
  );
  Adder m_353 ( // @[MUL.scala 102:19]
    .io_x1(m_353_io_x1),
    .io_x2(m_353_io_x2),
    .io_x3(m_353_io_x3),
    .io_s(m_353_io_s),
    .io_cout(m_353_io_cout)
  );
  Half_Adder m_354 ( // @[MUL.scala 124:19]
    .io_in_0(m_354_io_in_0),
    .io_in_1(m_354_io_in_1),
    .io_out_0(m_354_io_out_0),
    .io_out_1(m_354_io_out_1)
  );
  Adder m_355 ( // @[MUL.scala 102:19]
    .io_x1(m_355_io_x1),
    .io_x2(m_355_io_x2),
    .io_x3(m_355_io_x3),
    .io_s(m_355_io_s),
    .io_cout(m_355_io_cout)
  );
  Adder m_356 ( // @[MUL.scala 102:19]
    .io_x1(m_356_io_x1),
    .io_x2(m_356_io_x2),
    .io_x3(m_356_io_x3),
    .io_s(m_356_io_s),
    .io_cout(m_356_io_cout)
  );
  Half_Adder m_357 ( // @[MUL.scala 124:19]
    .io_in_0(m_357_io_in_0),
    .io_in_1(m_357_io_in_1),
    .io_out_0(m_357_io_out_0),
    .io_out_1(m_357_io_out_1)
  );
  Adder m_358 ( // @[MUL.scala 102:19]
    .io_x1(m_358_io_x1),
    .io_x2(m_358_io_x2),
    .io_x3(m_358_io_x3),
    .io_s(m_358_io_s),
    .io_cout(m_358_io_cout)
  );
  Adder m_359 ( // @[MUL.scala 102:19]
    .io_x1(m_359_io_x1),
    .io_x2(m_359_io_x2),
    .io_x3(m_359_io_x3),
    .io_s(m_359_io_s),
    .io_cout(m_359_io_cout)
  );
  Half_Adder m_360 ( // @[MUL.scala 124:19]
    .io_in_0(m_360_io_in_0),
    .io_in_1(m_360_io_in_1),
    .io_out_0(m_360_io_out_0),
    .io_out_1(m_360_io_out_1)
  );
  Adder m_361 ( // @[MUL.scala 102:19]
    .io_x1(m_361_io_x1),
    .io_x2(m_361_io_x2),
    .io_x3(m_361_io_x3),
    .io_s(m_361_io_s),
    .io_cout(m_361_io_cout)
  );
  Adder m_362 ( // @[MUL.scala 102:19]
    .io_x1(m_362_io_x1),
    .io_x2(m_362_io_x2),
    .io_x3(m_362_io_x3),
    .io_s(m_362_io_s),
    .io_cout(m_362_io_cout)
  );
  Adder m_363 ( // @[MUL.scala 102:19]
    .io_x1(m_363_io_x1),
    .io_x2(m_363_io_x2),
    .io_x3(m_363_io_x3),
    .io_s(m_363_io_s),
    .io_cout(m_363_io_cout)
  );
  Adder m_364 ( // @[MUL.scala 102:19]
    .io_x1(m_364_io_x1),
    .io_x2(m_364_io_x2),
    .io_x3(m_364_io_x3),
    .io_s(m_364_io_s),
    .io_cout(m_364_io_cout)
  );
  Adder m_365 ( // @[MUL.scala 102:19]
    .io_x1(m_365_io_x1),
    .io_x2(m_365_io_x2),
    .io_x3(m_365_io_x3),
    .io_s(m_365_io_s),
    .io_cout(m_365_io_cout)
  );
  Adder m_366 ( // @[MUL.scala 102:19]
    .io_x1(m_366_io_x1),
    .io_x2(m_366_io_x2),
    .io_x3(m_366_io_x3),
    .io_s(m_366_io_s),
    .io_cout(m_366_io_cout)
  );
  Adder m_367 ( // @[MUL.scala 102:19]
    .io_x1(m_367_io_x1),
    .io_x2(m_367_io_x2),
    .io_x3(m_367_io_x3),
    .io_s(m_367_io_s),
    .io_cout(m_367_io_cout)
  );
  Adder m_368 ( // @[MUL.scala 102:19]
    .io_x1(m_368_io_x1),
    .io_x2(m_368_io_x2),
    .io_x3(m_368_io_x3),
    .io_s(m_368_io_s),
    .io_cout(m_368_io_cout)
  );
  Adder m_369 ( // @[MUL.scala 102:19]
    .io_x1(m_369_io_x1),
    .io_x2(m_369_io_x2),
    .io_x3(m_369_io_x3),
    .io_s(m_369_io_s),
    .io_cout(m_369_io_cout)
  );
  Adder m_370 ( // @[MUL.scala 102:19]
    .io_x1(m_370_io_x1),
    .io_x2(m_370_io_x2),
    .io_x3(m_370_io_x3),
    .io_s(m_370_io_s),
    .io_cout(m_370_io_cout)
  );
  Adder m_371 ( // @[MUL.scala 102:19]
    .io_x1(m_371_io_x1),
    .io_x2(m_371_io_x2),
    .io_x3(m_371_io_x3),
    .io_s(m_371_io_s),
    .io_cout(m_371_io_cout)
  );
  Adder m_372 ( // @[MUL.scala 102:19]
    .io_x1(m_372_io_x1),
    .io_x2(m_372_io_x2),
    .io_x3(m_372_io_x3),
    .io_s(m_372_io_s),
    .io_cout(m_372_io_cout)
  );
  Adder m_373 ( // @[MUL.scala 102:19]
    .io_x1(m_373_io_x1),
    .io_x2(m_373_io_x2),
    .io_x3(m_373_io_x3),
    .io_s(m_373_io_s),
    .io_cout(m_373_io_cout)
  );
  Half_Adder m_374 ( // @[MUL.scala 124:19]
    .io_in_0(m_374_io_in_0),
    .io_in_1(m_374_io_in_1),
    .io_out_0(m_374_io_out_0),
    .io_out_1(m_374_io_out_1)
  );
  Adder m_375 ( // @[MUL.scala 102:19]
    .io_x1(m_375_io_x1),
    .io_x2(m_375_io_x2),
    .io_x3(m_375_io_x3),
    .io_s(m_375_io_s),
    .io_cout(m_375_io_cout)
  );
  Adder m_376 ( // @[MUL.scala 102:19]
    .io_x1(m_376_io_x1),
    .io_x2(m_376_io_x2),
    .io_x3(m_376_io_x3),
    .io_s(m_376_io_s),
    .io_cout(m_376_io_cout)
  );
  Adder m_377 ( // @[MUL.scala 102:19]
    .io_x1(m_377_io_x1),
    .io_x2(m_377_io_x2),
    .io_x3(m_377_io_x3),
    .io_s(m_377_io_s),
    .io_cout(m_377_io_cout)
  );
  Adder m_378 ( // @[MUL.scala 102:19]
    .io_x1(m_378_io_x1),
    .io_x2(m_378_io_x2),
    .io_x3(m_378_io_x3),
    .io_s(m_378_io_s),
    .io_cout(m_378_io_cout)
  );
  Adder m_379 ( // @[MUL.scala 102:19]
    .io_x1(m_379_io_x1),
    .io_x2(m_379_io_x2),
    .io_x3(m_379_io_x3),
    .io_s(m_379_io_s),
    .io_cout(m_379_io_cout)
  );
  Adder m_380 ( // @[MUL.scala 102:19]
    .io_x1(m_380_io_x1),
    .io_x2(m_380_io_x2),
    .io_x3(m_380_io_x3),
    .io_s(m_380_io_s),
    .io_cout(m_380_io_cout)
  );
  Half_Adder m_381 ( // @[MUL.scala 124:19]
    .io_in_0(m_381_io_in_0),
    .io_in_1(m_381_io_in_1),
    .io_out_0(m_381_io_out_0),
    .io_out_1(m_381_io_out_1)
  );
  Half_Adder m_382 ( // @[MUL.scala 124:19]
    .io_in_0(m_382_io_in_0),
    .io_in_1(m_382_io_in_1),
    .io_out_0(m_382_io_out_0),
    .io_out_1(m_382_io_out_1)
  );
  Half_Adder m_383 ( // @[MUL.scala 124:19]
    .io_in_0(m_383_io_in_0),
    .io_in_1(m_383_io_in_1),
    .io_out_0(m_383_io_out_0),
    .io_out_1(m_383_io_out_1)
  );
  Half_Adder m_384 ( // @[MUL.scala 124:19]
    .io_in_0(m_384_io_in_0),
    .io_in_1(m_384_io_in_1),
    .io_out_0(m_384_io_out_0),
    .io_out_1(m_384_io_out_1)
  );
  Half_Adder m_385 ( // @[MUL.scala 124:19]
    .io_in_0(m_385_io_in_0),
    .io_in_1(m_385_io_in_1),
    .io_out_0(m_385_io_out_0),
    .io_out_1(m_385_io_out_1)
  );
  Half_Adder m_386 ( // @[MUL.scala 124:19]
    .io_in_0(m_386_io_in_0),
    .io_in_1(m_386_io_in_1),
    .io_out_0(m_386_io_out_0),
    .io_out_1(m_386_io_out_1)
  );
  Half_Adder m_387 ( // @[MUL.scala 124:19]
    .io_in_0(m_387_io_in_0),
    .io_in_1(m_387_io_in_1),
    .io_out_0(m_387_io_out_0),
    .io_out_1(m_387_io_out_1)
  );
  Half_Adder m_388 ( // @[MUL.scala 124:19]
    .io_in_0(m_388_io_in_0),
    .io_in_1(m_388_io_in_1),
    .io_out_0(m_388_io_out_0),
    .io_out_1(m_388_io_out_1)
  );
  Half_Adder m_389 ( // @[MUL.scala 124:19]
    .io_in_0(m_389_io_in_0),
    .io_in_1(m_389_io_in_1),
    .io_out_0(m_389_io_out_0),
    .io_out_1(m_389_io_out_1)
  );
  Half_Adder m_390 ( // @[MUL.scala 124:19]
    .io_in_0(m_390_io_in_0),
    .io_in_1(m_390_io_in_1),
    .io_out_0(m_390_io_out_0),
    .io_out_1(m_390_io_out_1)
  );
  Adder m_391 ( // @[MUL.scala 102:19]
    .io_x1(m_391_io_x1),
    .io_x2(m_391_io_x2),
    .io_x3(m_391_io_x3),
    .io_s(m_391_io_s),
    .io_cout(m_391_io_cout)
  );
  Adder m_392 ( // @[MUL.scala 102:19]
    .io_x1(m_392_io_x1),
    .io_x2(m_392_io_x2),
    .io_x3(m_392_io_x3),
    .io_s(m_392_io_s),
    .io_cout(m_392_io_cout)
  );
  Adder m_393 ( // @[MUL.scala 102:19]
    .io_x1(m_393_io_x1),
    .io_x2(m_393_io_x2),
    .io_x3(m_393_io_x3),
    .io_s(m_393_io_s),
    .io_cout(m_393_io_cout)
  );
  Adder m_394 ( // @[MUL.scala 102:19]
    .io_x1(m_394_io_x1),
    .io_x2(m_394_io_x2),
    .io_x3(m_394_io_x3),
    .io_s(m_394_io_s),
    .io_cout(m_394_io_cout)
  );
  Adder m_395 ( // @[MUL.scala 102:19]
    .io_x1(m_395_io_x1),
    .io_x2(m_395_io_x2),
    .io_x3(m_395_io_x3),
    .io_s(m_395_io_s),
    .io_cout(m_395_io_cout)
  );
  Adder m_396 ( // @[MUL.scala 102:19]
    .io_x1(m_396_io_x1),
    .io_x2(m_396_io_x2),
    .io_x3(m_396_io_x3),
    .io_s(m_396_io_s),
    .io_cout(m_396_io_cout)
  );
  Adder m_397 ( // @[MUL.scala 102:19]
    .io_x1(m_397_io_x1),
    .io_x2(m_397_io_x2),
    .io_x3(m_397_io_x3),
    .io_s(m_397_io_s),
    .io_cout(m_397_io_cout)
  );
  Adder m_398 ( // @[MUL.scala 102:19]
    .io_x1(m_398_io_x1),
    .io_x2(m_398_io_x2),
    .io_x3(m_398_io_x3),
    .io_s(m_398_io_s),
    .io_cout(m_398_io_cout)
  );
  Adder m_399 ( // @[MUL.scala 102:19]
    .io_x1(m_399_io_x1),
    .io_x2(m_399_io_x2),
    .io_x3(m_399_io_x3),
    .io_s(m_399_io_s),
    .io_cout(m_399_io_cout)
  );
  Adder m_400 ( // @[MUL.scala 102:19]
    .io_x1(m_400_io_x1),
    .io_x2(m_400_io_x2),
    .io_x3(m_400_io_x3),
    .io_s(m_400_io_s),
    .io_cout(m_400_io_cout)
  );
  Half_Adder m_401 ( // @[MUL.scala 124:19]
    .io_in_0(m_401_io_in_0),
    .io_in_1(m_401_io_in_1),
    .io_out_0(m_401_io_out_0),
    .io_out_1(m_401_io_out_1)
  );
  Adder m_402 ( // @[MUL.scala 102:19]
    .io_x1(m_402_io_x1),
    .io_x2(m_402_io_x2),
    .io_x3(m_402_io_x3),
    .io_s(m_402_io_s),
    .io_cout(m_402_io_cout)
  );
  Half_Adder m_403 ( // @[MUL.scala 124:19]
    .io_in_0(m_403_io_in_0),
    .io_in_1(m_403_io_in_1),
    .io_out_0(m_403_io_out_0),
    .io_out_1(m_403_io_out_1)
  );
  Adder m_404 ( // @[MUL.scala 102:19]
    .io_x1(m_404_io_x1),
    .io_x2(m_404_io_x2),
    .io_x3(m_404_io_x3),
    .io_s(m_404_io_s),
    .io_cout(m_404_io_cout)
  );
  Half_Adder m_405 ( // @[MUL.scala 124:19]
    .io_in_0(m_405_io_in_0),
    .io_in_1(m_405_io_in_1),
    .io_out_0(m_405_io_out_0),
    .io_out_1(m_405_io_out_1)
  );
  Adder m_406 ( // @[MUL.scala 102:19]
    .io_x1(m_406_io_x1),
    .io_x2(m_406_io_x2),
    .io_x3(m_406_io_x3),
    .io_s(m_406_io_s),
    .io_cout(m_406_io_cout)
  );
  Half_Adder m_407 ( // @[MUL.scala 124:19]
    .io_in_0(m_407_io_in_0),
    .io_in_1(m_407_io_in_1),
    .io_out_0(m_407_io_out_0),
    .io_out_1(m_407_io_out_1)
  );
  Adder m_408 ( // @[MUL.scala 102:19]
    .io_x1(m_408_io_x1),
    .io_x2(m_408_io_x2),
    .io_x3(m_408_io_x3),
    .io_s(m_408_io_s),
    .io_cout(m_408_io_cout)
  );
  Adder m_409 ( // @[MUL.scala 102:19]
    .io_x1(m_409_io_x1),
    .io_x2(m_409_io_x2),
    .io_x3(m_409_io_x3),
    .io_s(m_409_io_s),
    .io_cout(m_409_io_cout)
  );
  Adder m_410 ( // @[MUL.scala 102:19]
    .io_x1(m_410_io_x1),
    .io_x2(m_410_io_x2),
    .io_x3(m_410_io_x3),
    .io_s(m_410_io_s),
    .io_cout(m_410_io_cout)
  );
  Adder m_411 ( // @[MUL.scala 102:19]
    .io_x1(m_411_io_x1),
    .io_x2(m_411_io_x2),
    .io_x3(m_411_io_x3),
    .io_s(m_411_io_s),
    .io_cout(m_411_io_cout)
  );
  Adder m_412 ( // @[MUL.scala 102:19]
    .io_x1(m_412_io_x1),
    .io_x2(m_412_io_x2),
    .io_x3(m_412_io_x3),
    .io_s(m_412_io_s),
    .io_cout(m_412_io_cout)
  );
  Adder m_413 ( // @[MUL.scala 102:19]
    .io_x1(m_413_io_x1),
    .io_x2(m_413_io_x2),
    .io_x3(m_413_io_x3),
    .io_s(m_413_io_s),
    .io_cout(m_413_io_cout)
  );
  Adder m_414 ( // @[MUL.scala 102:19]
    .io_x1(m_414_io_x1),
    .io_x2(m_414_io_x2),
    .io_x3(m_414_io_x3),
    .io_s(m_414_io_s),
    .io_cout(m_414_io_cout)
  );
  Adder m_415 ( // @[MUL.scala 102:19]
    .io_x1(m_415_io_x1),
    .io_x2(m_415_io_x2),
    .io_x3(m_415_io_x3),
    .io_s(m_415_io_s),
    .io_cout(m_415_io_cout)
  );
  Adder m_416 ( // @[MUL.scala 102:19]
    .io_x1(m_416_io_x1),
    .io_x2(m_416_io_x2),
    .io_x3(m_416_io_x3),
    .io_s(m_416_io_s),
    .io_cout(m_416_io_cout)
  );
  Adder m_417 ( // @[MUL.scala 102:19]
    .io_x1(m_417_io_x1),
    .io_x2(m_417_io_x2),
    .io_x3(m_417_io_x3),
    .io_s(m_417_io_s),
    .io_cout(m_417_io_cout)
  );
  Adder m_418 ( // @[MUL.scala 102:19]
    .io_x1(m_418_io_x1),
    .io_x2(m_418_io_x2),
    .io_x3(m_418_io_x3),
    .io_s(m_418_io_s),
    .io_cout(m_418_io_cout)
  );
  Adder m_419 ( // @[MUL.scala 102:19]
    .io_x1(m_419_io_x1),
    .io_x2(m_419_io_x2),
    .io_x3(m_419_io_x3),
    .io_s(m_419_io_s),
    .io_cout(m_419_io_cout)
  );
  Adder m_420 ( // @[MUL.scala 102:19]
    .io_x1(m_420_io_x1),
    .io_x2(m_420_io_x2),
    .io_x3(m_420_io_x3),
    .io_s(m_420_io_s),
    .io_cout(m_420_io_cout)
  );
  Adder m_421 ( // @[MUL.scala 102:19]
    .io_x1(m_421_io_x1),
    .io_x2(m_421_io_x2),
    .io_x3(m_421_io_x3),
    .io_s(m_421_io_s),
    .io_cout(m_421_io_cout)
  );
  Adder m_422 ( // @[MUL.scala 102:19]
    .io_x1(m_422_io_x1),
    .io_x2(m_422_io_x2),
    .io_x3(m_422_io_x3),
    .io_s(m_422_io_s),
    .io_cout(m_422_io_cout)
  );
  Adder m_423 ( // @[MUL.scala 102:19]
    .io_x1(m_423_io_x1),
    .io_x2(m_423_io_x2),
    .io_x3(m_423_io_x3),
    .io_s(m_423_io_s),
    .io_cout(m_423_io_cout)
  );
  Adder m_424 ( // @[MUL.scala 102:19]
    .io_x1(m_424_io_x1),
    .io_x2(m_424_io_x2),
    .io_x3(m_424_io_x3),
    .io_s(m_424_io_s),
    .io_cout(m_424_io_cout)
  );
  Adder m_425 ( // @[MUL.scala 102:19]
    .io_x1(m_425_io_x1),
    .io_x2(m_425_io_x2),
    .io_x3(m_425_io_x3),
    .io_s(m_425_io_s),
    .io_cout(m_425_io_cout)
  );
  Adder m_426 ( // @[MUL.scala 102:19]
    .io_x1(m_426_io_x1),
    .io_x2(m_426_io_x2),
    .io_x3(m_426_io_x3),
    .io_s(m_426_io_s),
    .io_cout(m_426_io_cout)
  );
  Adder m_427 ( // @[MUL.scala 102:19]
    .io_x1(m_427_io_x1),
    .io_x2(m_427_io_x2),
    .io_x3(m_427_io_x3),
    .io_s(m_427_io_s),
    .io_cout(m_427_io_cout)
  );
  Half_Adder m_428 ( // @[MUL.scala 124:19]
    .io_in_0(m_428_io_in_0),
    .io_in_1(m_428_io_in_1),
    .io_out_0(m_428_io_out_0),
    .io_out_1(m_428_io_out_1)
  );
  Adder m_429 ( // @[MUL.scala 102:19]
    .io_x1(m_429_io_x1),
    .io_x2(m_429_io_x2),
    .io_x3(m_429_io_x3),
    .io_s(m_429_io_s),
    .io_cout(m_429_io_cout)
  );
  Adder m_430 ( // @[MUL.scala 102:19]
    .io_x1(m_430_io_x1),
    .io_x2(m_430_io_x2),
    .io_x3(m_430_io_x3),
    .io_s(m_430_io_s),
    .io_cout(m_430_io_cout)
  );
  Half_Adder m_431 ( // @[MUL.scala 124:19]
    .io_in_0(m_431_io_in_0),
    .io_in_1(m_431_io_in_1),
    .io_out_0(m_431_io_out_0),
    .io_out_1(m_431_io_out_1)
  );
  Adder m_432 ( // @[MUL.scala 102:19]
    .io_x1(m_432_io_x1),
    .io_x2(m_432_io_x2),
    .io_x3(m_432_io_x3),
    .io_s(m_432_io_s),
    .io_cout(m_432_io_cout)
  );
  Adder m_433 ( // @[MUL.scala 102:19]
    .io_x1(m_433_io_x1),
    .io_x2(m_433_io_x2),
    .io_x3(m_433_io_x3),
    .io_s(m_433_io_s),
    .io_cout(m_433_io_cout)
  );
  Half_Adder m_434 ( // @[MUL.scala 124:19]
    .io_in_0(m_434_io_in_0),
    .io_in_1(m_434_io_in_1),
    .io_out_0(m_434_io_out_0),
    .io_out_1(m_434_io_out_1)
  );
  Adder m_435 ( // @[MUL.scala 102:19]
    .io_x1(m_435_io_x1),
    .io_x2(m_435_io_x2),
    .io_x3(m_435_io_x3),
    .io_s(m_435_io_s),
    .io_cout(m_435_io_cout)
  );
  Adder m_436 ( // @[MUL.scala 102:19]
    .io_x1(m_436_io_x1),
    .io_x2(m_436_io_x2),
    .io_x3(m_436_io_x3),
    .io_s(m_436_io_s),
    .io_cout(m_436_io_cout)
  );
  Half_Adder m_437 ( // @[MUL.scala 124:19]
    .io_in_0(m_437_io_in_0),
    .io_in_1(m_437_io_in_1),
    .io_out_0(m_437_io_out_0),
    .io_out_1(m_437_io_out_1)
  );
  Adder m_438 ( // @[MUL.scala 102:19]
    .io_x1(m_438_io_x1),
    .io_x2(m_438_io_x2),
    .io_x3(m_438_io_x3),
    .io_s(m_438_io_s),
    .io_cout(m_438_io_cout)
  );
  Adder m_439 ( // @[MUL.scala 102:19]
    .io_x1(m_439_io_x1),
    .io_x2(m_439_io_x2),
    .io_x3(m_439_io_x3),
    .io_s(m_439_io_s),
    .io_cout(m_439_io_cout)
  );
  Half_Adder m_440 ( // @[MUL.scala 124:19]
    .io_in_0(m_440_io_in_0),
    .io_in_1(m_440_io_in_1),
    .io_out_0(m_440_io_out_0),
    .io_out_1(m_440_io_out_1)
  );
  Adder m_441 ( // @[MUL.scala 102:19]
    .io_x1(m_441_io_x1),
    .io_x2(m_441_io_x2),
    .io_x3(m_441_io_x3),
    .io_s(m_441_io_s),
    .io_cout(m_441_io_cout)
  );
  Adder m_442 ( // @[MUL.scala 102:19]
    .io_x1(m_442_io_x1),
    .io_x2(m_442_io_x2),
    .io_x3(m_442_io_x3),
    .io_s(m_442_io_s),
    .io_cout(m_442_io_cout)
  );
  Half_Adder m_443 ( // @[MUL.scala 124:19]
    .io_in_0(m_443_io_in_0),
    .io_in_1(m_443_io_in_1),
    .io_out_0(m_443_io_out_0),
    .io_out_1(m_443_io_out_1)
  );
  Adder m_444 ( // @[MUL.scala 102:19]
    .io_x1(m_444_io_x1),
    .io_x2(m_444_io_x2),
    .io_x3(m_444_io_x3),
    .io_s(m_444_io_s),
    .io_cout(m_444_io_cout)
  );
  Adder m_445 ( // @[MUL.scala 102:19]
    .io_x1(m_445_io_x1),
    .io_x2(m_445_io_x2),
    .io_x3(m_445_io_x3),
    .io_s(m_445_io_s),
    .io_cout(m_445_io_cout)
  );
  Half_Adder m_446 ( // @[MUL.scala 124:19]
    .io_in_0(m_446_io_in_0),
    .io_in_1(m_446_io_in_1),
    .io_out_0(m_446_io_out_0),
    .io_out_1(m_446_io_out_1)
  );
  Adder m_447 ( // @[MUL.scala 102:19]
    .io_x1(m_447_io_x1),
    .io_x2(m_447_io_x2),
    .io_x3(m_447_io_x3),
    .io_s(m_447_io_s),
    .io_cout(m_447_io_cout)
  );
  Adder m_448 ( // @[MUL.scala 102:19]
    .io_x1(m_448_io_x1),
    .io_x2(m_448_io_x2),
    .io_x3(m_448_io_x3),
    .io_s(m_448_io_s),
    .io_cout(m_448_io_cout)
  );
  Half_Adder m_449 ( // @[MUL.scala 124:19]
    .io_in_0(m_449_io_in_0),
    .io_in_1(m_449_io_in_1),
    .io_out_0(m_449_io_out_0),
    .io_out_1(m_449_io_out_1)
  );
  Adder m_450 ( // @[MUL.scala 102:19]
    .io_x1(m_450_io_x1),
    .io_x2(m_450_io_x2),
    .io_x3(m_450_io_x3),
    .io_s(m_450_io_s),
    .io_cout(m_450_io_cout)
  );
  Adder m_451 ( // @[MUL.scala 102:19]
    .io_x1(m_451_io_x1),
    .io_x2(m_451_io_x2),
    .io_x3(m_451_io_x3),
    .io_s(m_451_io_s),
    .io_cout(m_451_io_cout)
  );
  Half_Adder m_452 ( // @[MUL.scala 124:19]
    .io_in_0(m_452_io_in_0),
    .io_in_1(m_452_io_in_1),
    .io_out_0(m_452_io_out_0),
    .io_out_1(m_452_io_out_1)
  );
  Adder m_453 ( // @[MUL.scala 102:19]
    .io_x1(m_453_io_x1),
    .io_x2(m_453_io_x2),
    .io_x3(m_453_io_x3),
    .io_s(m_453_io_s),
    .io_cout(m_453_io_cout)
  );
  Adder m_454 ( // @[MUL.scala 102:19]
    .io_x1(m_454_io_x1),
    .io_x2(m_454_io_x2),
    .io_x3(m_454_io_x3),
    .io_s(m_454_io_s),
    .io_cout(m_454_io_cout)
  );
  Half_Adder m_455 ( // @[MUL.scala 124:19]
    .io_in_0(m_455_io_in_0),
    .io_in_1(m_455_io_in_1),
    .io_out_0(m_455_io_out_0),
    .io_out_1(m_455_io_out_1)
  );
  Adder m_456 ( // @[MUL.scala 102:19]
    .io_x1(m_456_io_x1),
    .io_x2(m_456_io_x2),
    .io_x3(m_456_io_x3),
    .io_s(m_456_io_s),
    .io_cout(m_456_io_cout)
  );
  Adder m_457 ( // @[MUL.scala 102:19]
    .io_x1(m_457_io_x1),
    .io_x2(m_457_io_x2),
    .io_x3(m_457_io_x3),
    .io_s(m_457_io_s),
    .io_cout(m_457_io_cout)
  );
  Adder m_458 ( // @[MUL.scala 102:19]
    .io_x1(m_458_io_x1),
    .io_x2(m_458_io_x2),
    .io_x3(m_458_io_x3),
    .io_s(m_458_io_s),
    .io_cout(m_458_io_cout)
  );
  Adder m_459 ( // @[MUL.scala 102:19]
    .io_x1(m_459_io_x1),
    .io_x2(m_459_io_x2),
    .io_x3(m_459_io_x3),
    .io_s(m_459_io_s),
    .io_cout(m_459_io_cout)
  );
  Adder m_460 ( // @[MUL.scala 102:19]
    .io_x1(m_460_io_x1),
    .io_x2(m_460_io_x2),
    .io_x3(m_460_io_x3),
    .io_s(m_460_io_s),
    .io_cout(m_460_io_cout)
  );
  Adder m_461 ( // @[MUL.scala 102:19]
    .io_x1(m_461_io_x1),
    .io_x2(m_461_io_x2),
    .io_x3(m_461_io_x3),
    .io_s(m_461_io_s),
    .io_cout(m_461_io_cout)
  );
  Adder m_462 ( // @[MUL.scala 102:19]
    .io_x1(m_462_io_x1),
    .io_x2(m_462_io_x2),
    .io_x3(m_462_io_x3),
    .io_s(m_462_io_s),
    .io_cout(m_462_io_cout)
  );
  Adder m_463 ( // @[MUL.scala 102:19]
    .io_x1(m_463_io_x1),
    .io_x2(m_463_io_x2),
    .io_x3(m_463_io_x3),
    .io_s(m_463_io_s),
    .io_cout(m_463_io_cout)
  );
  Adder m_464 ( // @[MUL.scala 102:19]
    .io_x1(m_464_io_x1),
    .io_x2(m_464_io_x2),
    .io_x3(m_464_io_x3),
    .io_s(m_464_io_s),
    .io_cout(m_464_io_cout)
  );
  Adder m_465 ( // @[MUL.scala 102:19]
    .io_x1(m_465_io_x1),
    .io_x2(m_465_io_x2),
    .io_x3(m_465_io_x3),
    .io_s(m_465_io_s),
    .io_cout(m_465_io_cout)
  );
  Adder m_466 ( // @[MUL.scala 102:19]
    .io_x1(m_466_io_x1),
    .io_x2(m_466_io_x2),
    .io_x3(m_466_io_x3),
    .io_s(m_466_io_s),
    .io_cout(m_466_io_cout)
  );
  Adder m_467 ( // @[MUL.scala 102:19]
    .io_x1(m_467_io_x1),
    .io_x2(m_467_io_x2),
    .io_x3(m_467_io_x3),
    .io_s(m_467_io_s),
    .io_cout(m_467_io_cout)
  );
  Adder m_468 ( // @[MUL.scala 102:19]
    .io_x1(m_468_io_x1),
    .io_x2(m_468_io_x2),
    .io_x3(m_468_io_x3),
    .io_s(m_468_io_s),
    .io_cout(m_468_io_cout)
  );
  Adder m_469 ( // @[MUL.scala 102:19]
    .io_x1(m_469_io_x1),
    .io_x2(m_469_io_x2),
    .io_x3(m_469_io_x3),
    .io_s(m_469_io_s),
    .io_cout(m_469_io_cout)
  );
  Adder m_470 ( // @[MUL.scala 102:19]
    .io_x1(m_470_io_x1),
    .io_x2(m_470_io_x2),
    .io_x3(m_470_io_x3),
    .io_s(m_470_io_s),
    .io_cout(m_470_io_cout)
  );
  Adder m_471 ( // @[MUL.scala 102:19]
    .io_x1(m_471_io_x1),
    .io_x2(m_471_io_x2),
    .io_x3(m_471_io_x3),
    .io_s(m_471_io_s),
    .io_cout(m_471_io_cout)
  );
  Adder m_472 ( // @[MUL.scala 102:19]
    .io_x1(m_472_io_x1),
    .io_x2(m_472_io_x2),
    .io_x3(m_472_io_x3),
    .io_s(m_472_io_s),
    .io_cout(m_472_io_cout)
  );
  Adder m_473 ( // @[MUL.scala 102:19]
    .io_x1(m_473_io_x1),
    .io_x2(m_473_io_x2),
    .io_x3(m_473_io_x3),
    .io_s(m_473_io_s),
    .io_cout(m_473_io_cout)
  );
  Adder m_474 ( // @[MUL.scala 102:19]
    .io_x1(m_474_io_x1),
    .io_x2(m_474_io_x2),
    .io_x3(m_474_io_x3),
    .io_s(m_474_io_s),
    .io_cout(m_474_io_cout)
  );
  Adder m_475 ( // @[MUL.scala 102:19]
    .io_x1(m_475_io_x1),
    .io_x2(m_475_io_x2),
    .io_x3(m_475_io_x3),
    .io_s(m_475_io_s),
    .io_cout(m_475_io_cout)
  );
  Adder m_476 ( // @[MUL.scala 102:19]
    .io_x1(m_476_io_x1),
    .io_x2(m_476_io_x2),
    .io_x3(m_476_io_x3),
    .io_s(m_476_io_s),
    .io_cout(m_476_io_cout)
  );
  Adder m_477 ( // @[MUL.scala 102:19]
    .io_x1(m_477_io_x1),
    .io_x2(m_477_io_x2),
    .io_x3(m_477_io_x3),
    .io_s(m_477_io_s),
    .io_cout(m_477_io_cout)
  );
  Adder m_478 ( // @[MUL.scala 102:19]
    .io_x1(m_478_io_x1),
    .io_x2(m_478_io_x2),
    .io_x3(m_478_io_x3),
    .io_s(m_478_io_s),
    .io_cout(m_478_io_cout)
  );
  Adder m_479 ( // @[MUL.scala 102:19]
    .io_x1(m_479_io_x1),
    .io_x2(m_479_io_x2),
    .io_x3(m_479_io_x3),
    .io_s(m_479_io_s),
    .io_cout(m_479_io_cout)
  );
  Adder m_480 ( // @[MUL.scala 102:19]
    .io_x1(m_480_io_x1),
    .io_x2(m_480_io_x2),
    .io_x3(m_480_io_x3),
    .io_s(m_480_io_s),
    .io_cout(m_480_io_cout)
  );
  Adder m_481 ( // @[MUL.scala 102:19]
    .io_x1(m_481_io_x1),
    .io_x2(m_481_io_x2),
    .io_x3(m_481_io_x3),
    .io_s(m_481_io_s),
    .io_cout(m_481_io_cout)
  );
  Adder m_482 ( // @[MUL.scala 102:19]
    .io_x1(m_482_io_x1),
    .io_x2(m_482_io_x2),
    .io_x3(m_482_io_x3),
    .io_s(m_482_io_s),
    .io_cout(m_482_io_cout)
  );
  Adder m_483 ( // @[MUL.scala 102:19]
    .io_x1(m_483_io_x1),
    .io_x2(m_483_io_x2),
    .io_x3(m_483_io_x3),
    .io_s(m_483_io_s),
    .io_cout(m_483_io_cout)
  );
  Adder m_484 ( // @[MUL.scala 102:19]
    .io_x1(m_484_io_x1),
    .io_x2(m_484_io_x2),
    .io_x3(m_484_io_x3),
    .io_s(m_484_io_s),
    .io_cout(m_484_io_cout)
  );
  Adder m_485 ( // @[MUL.scala 102:19]
    .io_x1(m_485_io_x1),
    .io_x2(m_485_io_x2),
    .io_x3(m_485_io_x3),
    .io_s(m_485_io_s),
    .io_cout(m_485_io_cout)
  );
  Adder m_486 ( // @[MUL.scala 102:19]
    .io_x1(m_486_io_x1),
    .io_x2(m_486_io_x2),
    .io_x3(m_486_io_x3),
    .io_s(m_486_io_s),
    .io_cout(m_486_io_cout)
  );
  Adder m_487 ( // @[MUL.scala 102:19]
    .io_x1(m_487_io_x1),
    .io_x2(m_487_io_x2),
    .io_x3(m_487_io_x3),
    .io_s(m_487_io_s),
    .io_cout(m_487_io_cout)
  );
  Adder m_488 ( // @[MUL.scala 102:19]
    .io_x1(m_488_io_x1),
    .io_x2(m_488_io_x2),
    .io_x3(m_488_io_x3),
    .io_s(m_488_io_s),
    .io_cout(m_488_io_cout)
  );
  Half_Adder m_489 ( // @[MUL.scala 124:19]
    .io_in_0(m_489_io_in_0),
    .io_in_1(m_489_io_in_1),
    .io_out_0(m_489_io_out_0),
    .io_out_1(m_489_io_out_1)
  );
  Half_Adder m_490 ( // @[MUL.scala 124:19]
    .io_in_0(m_490_io_in_0),
    .io_in_1(m_490_io_in_1),
    .io_out_0(m_490_io_out_0),
    .io_out_1(m_490_io_out_1)
  );
  Half_Adder m_491 ( // @[MUL.scala 124:19]
    .io_in_0(m_491_io_in_0),
    .io_in_1(m_491_io_in_1),
    .io_out_0(m_491_io_out_0),
    .io_out_1(m_491_io_out_1)
  );
  Half_Adder m_492 ( // @[MUL.scala 124:19]
    .io_in_0(m_492_io_in_0),
    .io_in_1(m_492_io_in_1),
    .io_out_0(m_492_io_out_0),
    .io_out_1(m_492_io_out_1)
  );
  Half_Adder m_493 ( // @[MUL.scala 124:19]
    .io_in_0(m_493_io_in_0),
    .io_in_1(m_493_io_in_1),
    .io_out_0(m_493_io_out_0),
    .io_out_1(m_493_io_out_1)
  );
  Half_Adder m_494 ( // @[MUL.scala 124:19]
    .io_in_0(m_494_io_in_0),
    .io_in_1(m_494_io_in_1),
    .io_out_0(m_494_io_out_0),
    .io_out_1(m_494_io_out_1)
  );
  Half_Adder m_495 ( // @[MUL.scala 124:19]
    .io_in_0(m_495_io_in_0),
    .io_in_1(m_495_io_in_1),
    .io_out_0(m_495_io_out_0),
    .io_out_1(m_495_io_out_1)
  );
  Half_Adder m_496 ( // @[MUL.scala 124:19]
    .io_in_0(m_496_io_in_0),
    .io_in_1(m_496_io_in_1),
    .io_out_0(m_496_io_out_0),
    .io_out_1(m_496_io_out_1)
  );
  Half_Adder m_497 ( // @[MUL.scala 124:19]
    .io_in_0(m_497_io_in_0),
    .io_in_1(m_497_io_in_1),
    .io_out_0(m_497_io_out_0),
    .io_out_1(m_497_io_out_1)
  );
  Half_Adder m_498 ( // @[MUL.scala 124:19]
    .io_in_0(m_498_io_in_0),
    .io_in_1(m_498_io_in_1),
    .io_out_0(m_498_io_out_0),
    .io_out_1(m_498_io_out_1)
  );
  Half_Adder m_499 ( // @[MUL.scala 124:19]
    .io_in_0(m_499_io_in_0),
    .io_in_1(m_499_io_in_1),
    .io_out_0(m_499_io_out_0),
    .io_out_1(m_499_io_out_1)
  );
  Half_Adder m_500 ( // @[MUL.scala 124:19]
    .io_in_0(m_500_io_in_0),
    .io_in_1(m_500_io_in_1),
    .io_out_0(m_500_io_out_0),
    .io_out_1(m_500_io_out_1)
  );
  Half_Adder m_501 ( // @[MUL.scala 124:19]
    .io_in_0(m_501_io_in_0),
    .io_in_1(m_501_io_in_1),
    .io_out_0(m_501_io_out_0),
    .io_out_1(m_501_io_out_1)
  );
  Half_Adder m_502 ( // @[MUL.scala 124:19]
    .io_in_0(m_502_io_in_0),
    .io_in_1(m_502_io_in_1),
    .io_out_0(m_502_io_out_0),
    .io_out_1(m_502_io_out_1)
  );
  Adder m_503 ( // @[MUL.scala 102:19]
    .io_x1(m_503_io_x1),
    .io_x2(m_503_io_x2),
    .io_x3(m_503_io_x3),
    .io_s(m_503_io_s),
    .io_cout(m_503_io_cout)
  );
  Adder m_504 ( // @[MUL.scala 102:19]
    .io_x1(m_504_io_x1),
    .io_x2(m_504_io_x2),
    .io_x3(m_504_io_x3),
    .io_s(m_504_io_s),
    .io_cout(m_504_io_cout)
  );
  Adder m_505 ( // @[MUL.scala 102:19]
    .io_x1(m_505_io_x1),
    .io_x2(m_505_io_x2),
    .io_x3(m_505_io_x3),
    .io_s(m_505_io_s),
    .io_cout(m_505_io_cout)
  );
  Adder m_506 ( // @[MUL.scala 102:19]
    .io_x1(m_506_io_x1),
    .io_x2(m_506_io_x2),
    .io_x3(m_506_io_x3),
    .io_s(m_506_io_s),
    .io_cout(m_506_io_cout)
  );
  Adder m_507 ( // @[MUL.scala 102:19]
    .io_x1(m_507_io_x1),
    .io_x2(m_507_io_x2),
    .io_x3(m_507_io_x3),
    .io_s(m_507_io_s),
    .io_cout(m_507_io_cout)
  );
  Adder m_508 ( // @[MUL.scala 102:19]
    .io_x1(m_508_io_x1),
    .io_x2(m_508_io_x2),
    .io_x3(m_508_io_x3),
    .io_s(m_508_io_s),
    .io_cout(m_508_io_cout)
  );
  Adder m_509 ( // @[MUL.scala 102:19]
    .io_x1(m_509_io_x1),
    .io_x2(m_509_io_x2),
    .io_x3(m_509_io_x3),
    .io_s(m_509_io_s),
    .io_cout(m_509_io_cout)
  );
  Adder m_510 ( // @[MUL.scala 102:19]
    .io_x1(m_510_io_x1),
    .io_x2(m_510_io_x2),
    .io_x3(m_510_io_x3),
    .io_s(m_510_io_s),
    .io_cout(m_510_io_cout)
  );
  Adder m_511 ( // @[MUL.scala 102:19]
    .io_x1(m_511_io_x1),
    .io_x2(m_511_io_x2),
    .io_x3(m_511_io_x3),
    .io_s(m_511_io_s),
    .io_cout(m_511_io_cout)
  );
  Adder m_512 ( // @[MUL.scala 102:19]
    .io_x1(m_512_io_x1),
    .io_x2(m_512_io_x2),
    .io_x3(m_512_io_x3),
    .io_s(m_512_io_s),
    .io_cout(m_512_io_cout)
  );
  Adder m_513 ( // @[MUL.scala 102:19]
    .io_x1(m_513_io_x1),
    .io_x2(m_513_io_x2),
    .io_x3(m_513_io_x3),
    .io_s(m_513_io_s),
    .io_cout(m_513_io_cout)
  );
  Adder m_514 ( // @[MUL.scala 102:19]
    .io_x1(m_514_io_x1),
    .io_x2(m_514_io_x2),
    .io_x3(m_514_io_x3),
    .io_s(m_514_io_s),
    .io_cout(m_514_io_cout)
  );
  Adder m_515 ( // @[MUL.scala 102:19]
    .io_x1(m_515_io_x1),
    .io_x2(m_515_io_x2),
    .io_x3(m_515_io_x3),
    .io_s(m_515_io_s),
    .io_cout(m_515_io_cout)
  );
  Adder m_516 ( // @[MUL.scala 102:19]
    .io_x1(m_516_io_x1),
    .io_x2(m_516_io_x2),
    .io_x3(m_516_io_x3),
    .io_s(m_516_io_s),
    .io_cout(m_516_io_cout)
  );
  Adder m_517 ( // @[MUL.scala 102:19]
    .io_x1(m_517_io_x1),
    .io_x2(m_517_io_x2),
    .io_x3(m_517_io_x3),
    .io_s(m_517_io_s),
    .io_cout(m_517_io_cout)
  );
  Half_Adder m_518 ( // @[MUL.scala 124:19]
    .io_in_0(m_518_io_in_0),
    .io_in_1(m_518_io_in_1),
    .io_out_0(m_518_io_out_0),
    .io_out_1(m_518_io_out_1)
  );
  Adder m_519 ( // @[MUL.scala 102:19]
    .io_x1(m_519_io_x1),
    .io_x2(m_519_io_x2),
    .io_x3(m_519_io_x3),
    .io_s(m_519_io_s),
    .io_cout(m_519_io_cout)
  );
  Half_Adder m_520 ( // @[MUL.scala 124:19]
    .io_in_0(m_520_io_in_0),
    .io_in_1(m_520_io_in_1),
    .io_out_0(m_520_io_out_0),
    .io_out_1(m_520_io_out_1)
  );
  Adder m_521 ( // @[MUL.scala 102:19]
    .io_x1(m_521_io_x1),
    .io_x2(m_521_io_x2),
    .io_x3(m_521_io_x3),
    .io_s(m_521_io_s),
    .io_cout(m_521_io_cout)
  );
  Half_Adder m_522 ( // @[MUL.scala 124:19]
    .io_in_0(m_522_io_in_0),
    .io_in_1(m_522_io_in_1),
    .io_out_0(m_522_io_out_0),
    .io_out_1(m_522_io_out_1)
  );
  Adder m_523 ( // @[MUL.scala 102:19]
    .io_x1(m_523_io_x1),
    .io_x2(m_523_io_x2),
    .io_x3(m_523_io_x3),
    .io_s(m_523_io_s),
    .io_cout(m_523_io_cout)
  );
  Half_Adder m_524 ( // @[MUL.scala 124:19]
    .io_in_0(m_524_io_in_0),
    .io_in_1(m_524_io_in_1),
    .io_out_0(m_524_io_out_0),
    .io_out_1(m_524_io_out_1)
  );
  Adder m_525 ( // @[MUL.scala 102:19]
    .io_x1(m_525_io_x1),
    .io_x2(m_525_io_x2),
    .io_x3(m_525_io_x3),
    .io_s(m_525_io_s),
    .io_cout(m_525_io_cout)
  );
  Half_Adder m_526 ( // @[MUL.scala 124:19]
    .io_in_0(m_526_io_in_0),
    .io_in_1(m_526_io_in_1),
    .io_out_0(m_526_io_out_0),
    .io_out_1(m_526_io_out_1)
  );
  Adder m_527 ( // @[MUL.scala 102:19]
    .io_x1(m_527_io_x1),
    .io_x2(m_527_io_x2),
    .io_x3(m_527_io_x3),
    .io_s(m_527_io_s),
    .io_cout(m_527_io_cout)
  );
  Adder m_528 ( // @[MUL.scala 102:19]
    .io_x1(m_528_io_x1),
    .io_x2(m_528_io_x2),
    .io_x3(m_528_io_x3),
    .io_s(m_528_io_s),
    .io_cout(m_528_io_cout)
  );
  Adder m_529 ( // @[MUL.scala 102:19]
    .io_x1(m_529_io_x1),
    .io_x2(m_529_io_x2),
    .io_x3(m_529_io_x3),
    .io_s(m_529_io_s),
    .io_cout(m_529_io_cout)
  );
  Adder m_530 ( // @[MUL.scala 102:19]
    .io_x1(m_530_io_x1),
    .io_x2(m_530_io_x2),
    .io_x3(m_530_io_x3),
    .io_s(m_530_io_s),
    .io_cout(m_530_io_cout)
  );
  Adder m_531 ( // @[MUL.scala 102:19]
    .io_x1(m_531_io_x1),
    .io_x2(m_531_io_x2),
    .io_x3(m_531_io_x3),
    .io_s(m_531_io_s),
    .io_cout(m_531_io_cout)
  );
  Adder m_532 ( // @[MUL.scala 102:19]
    .io_x1(m_532_io_x1),
    .io_x2(m_532_io_x2),
    .io_x3(m_532_io_x3),
    .io_s(m_532_io_s),
    .io_cout(m_532_io_cout)
  );
  Adder m_533 ( // @[MUL.scala 102:19]
    .io_x1(m_533_io_x1),
    .io_x2(m_533_io_x2),
    .io_x3(m_533_io_x3),
    .io_s(m_533_io_s),
    .io_cout(m_533_io_cout)
  );
  Adder m_534 ( // @[MUL.scala 102:19]
    .io_x1(m_534_io_x1),
    .io_x2(m_534_io_x2),
    .io_x3(m_534_io_x3),
    .io_s(m_534_io_s),
    .io_cout(m_534_io_cout)
  );
  Adder m_535 ( // @[MUL.scala 102:19]
    .io_x1(m_535_io_x1),
    .io_x2(m_535_io_x2),
    .io_x3(m_535_io_x3),
    .io_s(m_535_io_s),
    .io_cout(m_535_io_cout)
  );
  Adder m_536 ( // @[MUL.scala 102:19]
    .io_x1(m_536_io_x1),
    .io_x2(m_536_io_x2),
    .io_x3(m_536_io_x3),
    .io_s(m_536_io_s),
    .io_cout(m_536_io_cout)
  );
  Adder m_537 ( // @[MUL.scala 102:19]
    .io_x1(m_537_io_x1),
    .io_x2(m_537_io_x2),
    .io_x3(m_537_io_x3),
    .io_s(m_537_io_s),
    .io_cout(m_537_io_cout)
  );
  Adder m_538 ( // @[MUL.scala 102:19]
    .io_x1(m_538_io_x1),
    .io_x2(m_538_io_x2),
    .io_x3(m_538_io_x3),
    .io_s(m_538_io_s),
    .io_cout(m_538_io_cout)
  );
  Adder m_539 ( // @[MUL.scala 102:19]
    .io_x1(m_539_io_x1),
    .io_x2(m_539_io_x2),
    .io_x3(m_539_io_x3),
    .io_s(m_539_io_s),
    .io_cout(m_539_io_cout)
  );
  Adder m_540 ( // @[MUL.scala 102:19]
    .io_x1(m_540_io_x1),
    .io_x2(m_540_io_x2),
    .io_x3(m_540_io_x3),
    .io_s(m_540_io_s),
    .io_cout(m_540_io_cout)
  );
  Adder m_541 ( // @[MUL.scala 102:19]
    .io_x1(m_541_io_x1),
    .io_x2(m_541_io_x2),
    .io_x3(m_541_io_x3),
    .io_s(m_541_io_s),
    .io_cout(m_541_io_cout)
  );
  Adder m_542 ( // @[MUL.scala 102:19]
    .io_x1(m_542_io_x1),
    .io_x2(m_542_io_x2),
    .io_x3(m_542_io_x3),
    .io_s(m_542_io_s),
    .io_cout(m_542_io_cout)
  );
  Adder m_543 ( // @[MUL.scala 102:19]
    .io_x1(m_543_io_x1),
    .io_x2(m_543_io_x2),
    .io_x3(m_543_io_x3),
    .io_s(m_543_io_s),
    .io_cout(m_543_io_cout)
  );
  Adder m_544 ( // @[MUL.scala 102:19]
    .io_x1(m_544_io_x1),
    .io_x2(m_544_io_x2),
    .io_x3(m_544_io_x3),
    .io_s(m_544_io_s),
    .io_cout(m_544_io_cout)
  );
  Adder m_545 ( // @[MUL.scala 102:19]
    .io_x1(m_545_io_x1),
    .io_x2(m_545_io_x2),
    .io_x3(m_545_io_x3),
    .io_s(m_545_io_s),
    .io_cout(m_545_io_cout)
  );
  Adder m_546 ( // @[MUL.scala 102:19]
    .io_x1(m_546_io_x1),
    .io_x2(m_546_io_x2),
    .io_x3(m_546_io_x3),
    .io_s(m_546_io_s),
    .io_cout(m_546_io_cout)
  );
  Adder m_547 ( // @[MUL.scala 102:19]
    .io_x1(m_547_io_x1),
    .io_x2(m_547_io_x2),
    .io_x3(m_547_io_x3),
    .io_s(m_547_io_s),
    .io_cout(m_547_io_cout)
  );
  Half_Adder m_548 ( // @[MUL.scala 124:19]
    .io_in_0(m_548_io_in_0),
    .io_in_1(m_548_io_in_1),
    .io_out_0(m_548_io_out_0),
    .io_out_1(m_548_io_out_1)
  );
  Adder m_549 ( // @[MUL.scala 102:19]
    .io_x1(m_549_io_x1),
    .io_x2(m_549_io_x2),
    .io_x3(m_549_io_x3),
    .io_s(m_549_io_s),
    .io_cout(m_549_io_cout)
  );
  Half_Adder m_550 ( // @[MUL.scala 124:19]
    .io_in_0(m_550_io_in_0),
    .io_in_1(m_550_io_in_1),
    .io_out_0(m_550_io_out_0),
    .io_out_1(m_550_io_out_1)
  );
  Adder m_551 ( // @[MUL.scala 102:19]
    .io_x1(m_551_io_x1),
    .io_x2(m_551_io_x2),
    .io_x3(m_551_io_x3),
    .io_s(m_551_io_s),
    .io_cout(m_551_io_cout)
  );
  Half_Adder m_552 ( // @[MUL.scala 124:19]
    .io_in_0(m_552_io_in_0),
    .io_in_1(m_552_io_in_1),
    .io_out_0(m_552_io_out_0),
    .io_out_1(m_552_io_out_1)
  );
  Adder m_553 ( // @[MUL.scala 102:19]
    .io_x1(m_553_io_x1),
    .io_x2(m_553_io_x2),
    .io_x3(m_553_io_x3),
    .io_s(m_553_io_s),
    .io_cout(m_553_io_cout)
  );
  Adder m_554 ( // @[MUL.scala 102:19]
    .io_x1(m_554_io_x1),
    .io_x2(m_554_io_x2),
    .io_x3(m_554_io_x3),
    .io_s(m_554_io_s),
    .io_cout(m_554_io_cout)
  );
  Adder m_555 ( // @[MUL.scala 102:19]
    .io_x1(m_555_io_x1),
    .io_x2(m_555_io_x2),
    .io_x3(m_555_io_x3),
    .io_s(m_555_io_s),
    .io_cout(m_555_io_cout)
  );
  Adder m_556 ( // @[MUL.scala 102:19]
    .io_x1(m_556_io_x1),
    .io_x2(m_556_io_x2),
    .io_x3(m_556_io_x3),
    .io_s(m_556_io_s),
    .io_cout(m_556_io_cout)
  );
  Adder m_557 ( // @[MUL.scala 102:19]
    .io_x1(m_557_io_x1),
    .io_x2(m_557_io_x2),
    .io_x3(m_557_io_x3),
    .io_s(m_557_io_s),
    .io_cout(m_557_io_cout)
  );
  Adder m_558 ( // @[MUL.scala 102:19]
    .io_x1(m_558_io_x1),
    .io_x2(m_558_io_x2),
    .io_x3(m_558_io_x3),
    .io_s(m_558_io_s),
    .io_cout(m_558_io_cout)
  );
  Adder m_559 ( // @[MUL.scala 102:19]
    .io_x1(m_559_io_x1),
    .io_x2(m_559_io_x2),
    .io_x3(m_559_io_x3),
    .io_s(m_559_io_s),
    .io_cout(m_559_io_cout)
  );
  Adder m_560 ( // @[MUL.scala 102:19]
    .io_x1(m_560_io_x1),
    .io_x2(m_560_io_x2),
    .io_x3(m_560_io_x3),
    .io_s(m_560_io_s),
    .io_cout(m_560_io_cout)
  );
  Adder m_561 ( // @[MUL.scala 102:19]
    .io_x1(m_561_io_x1),
    .io_x2(m_561_io_x2),
    .io_x3(m_561_io_x3),
    .io_s(m_561_io_s),
    .io_cout(m_561_io_cout)
  );
  Adder m_562 ( // @[MUL.scala 102:19]
    .io_x1(m_562_io_x1),
    .io_x2(m_562_io_x2),
    .io_x3(m_562_io_x3),
    .io_s(m_562_io_s),
    .io_cout(m_562_io_cout)
  );
  Adder m_563 ( // @[MUL.scala 102:19]
    .io_x1(m_563_io_x1),
    .io_x2(m_563_io_x2),
    .io_x3(m_563_io_x3),
    .io_s(m_563_io_s),
    .io_cout(m_563_io_cout)
  );
  Adder m_564 ( // @[MUL.scala 102:19]
    .io_x1(m_564_io_x1),
    .io_x2(m_564_io_x2),
    .io_x3(m_564_io_x3),
    .io_s(m_564_io_s),
    .io_cout(m_564_io_cout)
  );
  Adder m_565 ( // @[MUL.scala 102:19]
    .io_x1(m_565_io_x1),
    .io_x2(m_565_io_x2),
    .io_x3(m_565_io_x3),
    .io_s(m_565_io_s),
    .io_cout(m_565_io_cout)
  );
  Adder m_566 ( // @[MUL.scala 102:19]
    .io_x1(m_566_io_x1),
    .io_x2(m_566_io_x2),
    .io_x3(m_566_io_x3),
    .io_s(m_566_io_s),
    .io_cout(m_566_io_cout)
  );
  Half_Adder m_567 ( // @[MUL.scala 124:19]
    .io_in_0(m_567_io_in_0),
    .io_in_1(m_567_io_in_1),
    .io_out_0(m_567_io_out_0),
    .io_out_1(m_567_io_out_1)
  );
  Half_Adder m_568 ( // @[MUL.scala 124:19]
    .io_in_0(m_568_io_in_0),
    .io_in_1(m_568_io_in_1),
    .io_out_0(m_568_io_out_0),
    .io_out_1(m_568_io_out_1)
  );
  Half_Adder m_569 ( // @[MUL.scala 124:19]
    .io_in_0(m_569_io_in_0),
    .io_in_1(m_569_io_in_1),
    .io_out_0(m_569_io_out_0),
    .io_out_1(m_569_io_out_1)
  );
  Half_Adder m_570 ( // @[MUL.scala 124:19]
    .io_in_0(m_570_io_in_0),
    .io_in_1(m_570_io_in_1),
    .io_out_0(m_570_io_out_0),
    .io_out_1(m_570_io_out_1)
  );
  Half_Adder m_571 ( // @[MUL.scala 124:19]
    .io_in_0(m_571_io_in_0),
    .io_in_1(m_571_io_in_1),
    .io_out_0(m_571_io_out_0),
    .io_out_1(m_571_io_out_1)
  );
  Half_Adder m_572 ( // @[MUL.scala 124:19]
    .io_in_0(m_572_io_in_0),
    .io_in_1(m_572_io_in_1),
    .io_out_0(m_572_io_out_0),
    .io_out_1(m_572_io_out_1)
  );
  Half_Adder m_573 ( // @[MUL.scala 124:19]
    .io_in_0(m_573_io_in_0),
    .io_in_1(m_573_io_in_1),
    .io_out_0(m_573_io_out_0),
    .io_out_1(m_573_io_out_1)
  );
  Half_Adder m_574 ( // @[MUL.scala 124:19]
    .io_in_0(m_574_io_in_0),
    .io_in_1(m_574_io_in_1),
    .io_out_0(m_574_io_out_0),
    .io_out_1(m_574_io_out_1)
  );
  Half_Adder m_575 ( // @[MUL.scala 124:19]
    .io_in_0(m_575_io_in_0),
    .io_in_1(m_575_io_in_1),
    .io_out_0(m_575_io_out_0),
    .io_out_1(m_575_io_out_1)
  );
  Half_Adder m_576 ( // @[MUL.scala 124:19]
    .io_in_0(m_576_io_in_0),
    .io_in_1(m_576_io_in_1),
    .io_out_0(m_576_io_out_0),
    .io_out_1(m_576_io_out_1)
  );
  Half_Adder m_577 ( // @[MUL.scala 124:19]
    .io_in_0(m_577_io_in_0),
    .io_in_1(m_577_io_in_1),
    .io_out_0(m_577_io_out_0),
    .io_out_1(m_577_io_out_1)
  );
  Half_Adder m_578 ( // @[MUL.scala 124:19]
    .io_in_0(m_578_io_in_0),
    .io_in_1(m_578_io_in_1),
    .io_out_0(m_578_io_out_0),
    .io_out_1(m_578_io_out_1)
  );
  Half_Adder m_579 ( // @[MUL.scala 124:19]
    .io_in_0(m_579_io_in_0),
    .io_in_1(m_579_io_in_1),
    .io_out_0(m_579_io_out_0),
    .io_out_1(m_579_io_out_1)
  );
  Half_Adder m_580 ( // @[MUL.scala 124:19]
    .io_in_0(m_580_io_in_0),
    .io_in_1(m_580_io_in_1),
    .io_out_0(m_580_io_out_0),
    .io_out_1(m_580_io_out_1)
  );
  Half_Adder m_581 ( // @[MUL.scala 124:19]
    .io_in_0(m_581_io_in_0),
    .io_in_1(m_581_io_in_1),
    .io_out_0(m_581_io_out_0),
    .io_out_1(m_581_io_out_1)
  );
  Half_Adder m_582 ( // @[MUL.scala 124:19]
    .io_in_0(m_582_io_in_0),
    .io_in_1(m_582_io_in_1),
    .io_out_0(m_582_io_out_0),
    .io_out_1(m_582_io_out_1)
  );
  Half_Adder m_583 ( // @[MUL.scala 124:19]
    .io_in_0(m_583_io_in_0),
    .io_in_1(m_583_io_in_1),
    .io_out_0(m_583_io_out_0),
    .io_out_1(m_583_io_out_1)
  );
  Half_Adder m_584 ( // @[MUL.scala 124:19]
    .io_in_0(m_584_io_in_0),
    .io_in_1(m_584_io_in_1),
    .io_out_0(m_584_io_out_0),
    .io_out_1(m_584_io_out_1)
  );
  Half_Adder m_585 ( // @[MUL.scala 124:19]
    .io_in_0(m_585_io_in_0),
    .io_in_1(m_585_io_in_1),
    .io_out_0(m_585_io_out_0),
    .io_out_1(m_585_io_out_1)
  );
  Half_Adder m_586 ( // @[MUL.scala 124:19]
    .io_in_0(m_586_io_in_0),
    .io_in_1(m_586_io_in_1),
    .io_out_0(m_586_io_out_0),
    .io_out_1(m_586_io_out_1)
  );
  Half_Adder m_587 ( // @[MUL.scala 124:19]
    .io_in_0(m_587_io_in_0),
    .io_in_1(m_587_io_in_1),
    .io_out_0(m_587_io_out_0),
    .io_out_1(m_587_io_out_1)
  );
  Half_Adder m_588 ( // @[MUL.scala 124:19]
    .io_in_0(m_588_io_in_0),
    .io_in_1(m_588_io_in_1),
    .io_out_0(m_588_io_out_0),
    .io_out_1(m_588_io_out_1)
  );
  Half_Adder m_589 ( // @[MUL.scala 124:19]
    .io_in_0(m_589_io_in_0),
    .io_in_1(m_589_io_in_1),
    .io_out_0(m_589_io_out_0),
    .io_out_1(m_589_io_out_1)
  );
  Adder m_590 ( // @[MUL.scala 102:19]
    .io_x1(m_590_io_x1),
    .io_x2(m_590_io_x2),
    .io_x3(m_590_io_x3),
    .io_s(m_590_io_s),
    .io_cout(m_590_io_cout)
  );
  Adder m_591 ( // @[MUL.scala 102:19]
    .io_x1(m_591_io_x1),
    .io_x2(m_591_io_x2),
    .io_x3(m_591_io_x3),
    .io_s(m_591_io_s),
    .io_cout(m_591_io_cout)
  );
  Adder m_592 ( // @[MUL.scala 102:19]
    .io_x1(m_592_io_x1),
    .io_x2(m_592_io_x2),
    .io_x3(m_592_io_x3),
    .io_s(m_592_io_s),
    .io_cout(m_592_io_cout)
  );
  Adder m_593 ( // @[MUL.scala 102:19]
    .io_x1(m_593_io_x1),
    .io_x2(m_593_io_x2),
    .io_x3(m_593_io_x3),
    .io_s(m_593_io_s),
    .io_cout(m_593_io_cout)
  );
  Adder m_594 ( // @[MUL.scala 102:19]
    .io_x1(m_594_io_x1),
    .io_x2(m_594_io_x2),
    .io_x3(m_594_io_x3),
    .io_s(m_594_io_s),
    .io_cout(m_594_io_cout)
  );
  Adder m_595 ( // @[MUL.scala 102:19]
    .io_x1(m_595_io_x1),
    .io_x2(m_595_io_x2),
    .io_x3(m_595_io_x3),
    .io_s(m_595_io_s),
    .io_cout(m_595_io_cout)
  );
  Adder m_596 ( // @[MUL.scala 102:19]
    .io_x1(m_596_io_x1),
    .io_x2(m_596_io_x2),
    .io_x3(m_596_io_x3),
    .io_s(m_596_io_s),
    .io_cout(m_596_io_cout)
  );
  Adder m_597 ( // @[MUL.scala 102:19]
    .io_x1(m_597_io_x1),
    .io_x2(m_597_io_x2),
    .io_x3(m_597_io_x3),
    .io_s(m_597_io_s),
    .io_cout(m_597_io_cout)
  );
  Adder m_598 ( // @[MUL.scala 102:19]
    .io_x1(m_598_io_x1),
    .io_x2(m_598_io_x2),
    .io_x3(m_598_io_x3),
    .io_s(m_598_io_s),
    .io_cout(m_598_io_cout)
  );
  Adder m_599 ( // @[MUL.scala 102:19]
    .io_x1(m_599_io_x1),
    .io_x2(m_599_io_x2),
    .io_x3(m_599_io_x3),
    .io_s(m_599_io_s),
    .io_cout(m_599_io_cout)
  );
  Adder m_600 ( // @[MUL.scala 102:19]
    .io_x1(m_600_io_x1),
    .io_x2(m_600_io_x2),
    .io_x3(m_600_io_x3),
    .io_s(m_600_io_s),
    .io_cout(m_600_io_cout)
  );
  Adder m_601 ( // @[MUL.scala 102:19]
    .io_x1(m_601_io_x1),
    .io_x2(m_601_io_x2),
    .io_x3(m_601_io_x3),
    .io_s(m_601_io_s),
    .io_cout(m_601_io_cout)
  );
  Adder m_602 ( // @[MUL.scala 102:19]
    .io_x1(m_602_io_x1),
    .io_x2(m_602_io_x2),
    .io_x3(m_602_io_x3),
    .io_s(m_602_io_s),
    .io_cout(m_602_io_cout)
  );
  Adder m_603 ( // @[MUL.scala 102:19]
    .io_x1(m_603_io_x1),
    .io_x2(m_603_io_x2),
    .io_x3(m_603_io_x3),
    .io_s(m_603_io_s),
    .io_cout(m_603_io_cout)
  );
  Adder m_604 ( // @[MUL.scala 102:19]
    .io_x1(m_604_io_x1),
    .io_x2(m_604_io_x2),
    .io_x3(m_604_io_x3),
    .io_s(m_604_io_s),
    .io_cout(m_604_io_cout)
  );
  Adder m_605 ( // @[MUL.scala 102:19]
    .io_x1(m_605_io_x1),
    .io_x2(m_605_io_x2),
    .io_x3(m_605_io_x3),
    .io_s(m_605_io_s),
    .io_cout(m_605_io_cout)
  );
  Adder m_606 ( // @[MUL.scala 102:19]
    .io_x1(m_606_io_x1),
    .io_x2(m_606_io_x2),
    .io_x3(m_606_io_x3),
    .io_s(m_606_io_s),
    .io_cout(m_606_io_cout)
  );
  Adder m_607 ( // @[MUL.scala 102:19]
    .io_x1(m_607_io_x1),
    .io_x2(m_607_io_x2),
    .io_x3(m_607_io_x3),
    .io_s(m_607_io_s),
    .io_cout(m_607_io_cout)
  );
  Adder m_608 ( // @[MUL.scala 102:19]
    .io_x1(m_608_io_x1),
    .io_x2(m_608_io_x2),
    .io_x3(m_608_io_x3),
    .io_s(m_608_io_s),
    .io_cout(m_608_io_cout)
  );
  Adder m_609 ( // @[MUL.scala 102:19]
    .io_x1(m_609_io_x1),
    .io_x2(m_609_io_x2),
    .io_x3(m_609_io_x3),
    .io_s(m_609_io_s),
    .io_cout(m_609_io_cout)
  );
  Adder m_610 ( // @[MUL.scala 102:19]
    .io_x1(m_610_io_x1),
    .io_x2(m_610_io_x2),
    .io_x3(m_610_io_x3),
    .io_s(m_610_io_s),
    .io_cout(m_610_io_cout)
  );
  Adder m_611 ( // @[MUL.scala 102:19]
    .io_x1(m_611_io_x1),
    .io_x2(m_611_io_x2),
    .io_x3(m_611_io_x3),
    .io_s(m_611_io_s),
    .io_cout(m_611_io_cout)
  );
  Adder m_612 ( // @[MUL.scala 102:19]
    .io_x1(m_612_io_x1),
    .io_x2(m_612_io_x2),
    .io_x3(m_612_io_x3),
    .io_s(m_612_io_s),
    .io_cout(m_612_io_cout)
  );
  Adder m_613 ( // @[MUL.scala 102:19]
    .io_x1(m_613_io_x1),
    .io_x2(m_613_io_x2),
    .io_x3(m_613_io_x3),
    .io_s(m_613_io_s),
    .io_cout(m_613_io_cout)
  );
  Adder m_614 ( // @[MUL.scala 102:19]
    .io_x1(m_614_io_x1),
    .io_x2(m_614_io_x2),
    .io_x3(m_614_io_x3),
    .io_s(m_614_io_s),
    .io_cout(m_614_io_cout)
  );
  Adder m_615 ( // @[MUL.scala 102:19]
    .io_x1(m_615_io_x1),
    .io_x2(m_615_io_x2),
    .io_x3(m_615_io_x3),
    .io_s(m_615_io_s),
    .io_cout(m_615_io_cout)
  );
  Adder m_616 ( // @[MUL.scala 102:19]
    .io_x1(m_616_io_x1),
    .io_x2(m_616_io_x2),
    .io_x3(m_616_io_x3),
    .io_s(m_616_io_s),
    .io_cout(m_616_io_cout)
  );
  Adder m_617 ( // @[MUL.scala 102:19]
    .io_x1(m_617_io_x1),
    .io_x2(m_617_io_x2),
    .io_x3(m_617_io_x3),
    .io_s(m_617_io_s),
    .io_cout(m_617_io_cout)
  );
  Adder m_618 ( // @[MUL.scala 102:19]
    .io_x1(m_618_io_x1),
    .io_x2(m_618_io_x2),
    .io_x3(m_618_io_x3),
    .io_s(m_618_io_s),
    .io_cout(m_618_io_cout)
  );
  Adder m_619 ( // @[MUL.scala 102:19]
    .io_x1(m_619_io_x1),
    .io_x2(m_619_io_x2),
    .io_x3(m_619_io_x3),
    .io_s(m_619_io_s),
    .io_cout(m_619_io_cout)
  );
  Adder m_620 ( // @[MUL.scala 102:19]
    .io_x1(m_620_io_x1),
    .io_x2(m_620_io_x2),
    .io_x3(m_620_io_x3),
    .io_s(m_620_io_s),
    .io_cout(m_620_io_cout)
  );
  Adder m_621 ( // @[MUL.scala 102:19]
    .io_x1(m_621_io_x1),
    .io_x2(m_621_io_x2),
    .io_x3(m_621_io_x3),
    .io_s(m_621_io_s),
    .io_cout(m_621_io_cout)
  );
  Adder m_622 ( // @[MUL.scala 102:19]
    .io_x1(m_622_io_x1),
    .io_x2(m_622_io_x2),
    .io_x3(m_622_io_x3),
    .io_s(m_622_io_s),
    .io_cout(m_622_io_cout)
  );
  Adder m_623 ( // @[MUL.scala 102:19]
    .io_x1(m_623_io_x1),
    .io_x2(m_623_io_x2),
    .io_x3(m_623_io_x3),
    .io_s(m_623_io_s),
    .io_cout(m_623_io_cout)
  );
  Half_Adder m_624 ( // @[MUL.scala 124:19]
    .io_in_0(m_624_io_in_0),
    .io_in_1(m_624_io_in_1),
    .io_out_0(m_624_io_out_0),
    .io_out_1(m_624_io_out_1)
  );
  Half_Adder m_625 ( // @[MUL.scala 124:19]
    .io_in_0(m_625_io_in_0),
    .io_in_1(m_625_io_in_1),
    .io_out_0(m_625_io_out_0),
    .io_out_1(m_625_io_out_1)
  );
  Half_Adder m_626 ( // @[MUL.scala 124:19]
    .io_in_0(m_626_io_in_0),
    .io_in_1(m_626_io_in_1),
    .io_out_0(m_626_io_out_0),
    .io_out_1(m_626_io_out_1)
  );
  Half_Adder m_627 ( // @[MUL.scala 124:19]
    .io_in_0(m_627_io_in_0),
    .io_in_1(m_627_io_in_1),
    .io_out_0(m_627_io_out_0),
    .io_out_1(m_627_io_out_1)
  );
  Half_Adder m_628 ( // @[MUL.scala 124:19]
    .io_in_0(m_628_io_in_0),
    .io_in_1(m_628_io_in_1),
    .io_out_0(m_628_io_out_0),
    .io_out_1(m_628_io_out_1)
  );
  Half_Adder m_629 ( // @[MUL.scala 124:19]
    .io_in_0(m_629_io_in_0),
    .io_in_1(m_629_io_in_1),
    .io_out_0(m_629_io_out_0),
    .io_out_1(m_629_io_out_1)
  );
  Half_Adder m_630 ( // @[MUL.scala 124:19]
    .io_in_0(m_630_io_in_0),
    .io_in_1(m_630_io_in_1),
    .io_out_0(m_630_io_out_0),
    .io_out_1(m_630_io_out_1)
  );
  Half_Adder m_631 ( // @[MUL.scala 124:19]
    .io_in_0(m_631_io_in_0),
    .io_in_1(m_631_io_in_1),
    .io_out_0(m_631_io_out_0),
    .io_out_1(m_631_io_out_1)
  );
  Half_Adder m_632 ( // @[MUL.scala 124:19]
    .io_in_0(m_632_io_in_0),
    .io_in_1(m_632_io_in_1),
    .io_out_0(m_632_io_out_0),
    .io_out_1(m_632_io_out_1)
  );
  Half_Adder m_633 ( // @[MUL.scala 124:19]
    .io_in_0(m_633_io_in_0),
    .io_in_1(m_633_io_in_1),
    .io_out_0(m_633_io_out_0),
    .io_out_1(m_633_io_out_1)
  );
  Half_Adder m_634 ( // @[MUL.scala 124:19]
    .io_in_0(m_634_io_in_0),
    .io_in_1(m_634_io_in_1),
    .io_out_0(m_634_io_out_0),
    .io_out_1(m_634_io_out_1)
  );
  Half_Adder m_635 ( // @[MUL.scala 124:19]
    .io_in_0(m_635_io_in_0),
    .io_in_1(m_635_io_in_1),
    .io_out_0(m_635_io_out_0),
    .io_out_1(m_635_io_out_1)
  );
  Half_Adder m_636 ( // @[MUL.scala 124:19]
    .io_in_0(m_636_io_in_0),
    .io_in_1(m_636_io_in_1),
    .io_out_0(m_636_io_out_0),
    .io_out_1(m_636_io_out_1)
  );
  Half_Adder m_637 ( // @[MUL.scala 124:19]
    .io_in_0(m_637_io_in_0),
    .io_in_1(m_637_io_in_1),
    .io_out_0(m_637_io_out_0),
    .io_out_1(m_637_io_out_1)
  );
  Half_Adder m_638 ( // @[MUL.scala 124:19]
    .io_in_0(m_638_io_in_0),
    .io_in_1(m_638_io_in_1),
    .io_out_0(m_638_io_out_0),
    .io_out_1(m_638_io_out_1)
  );
  Half_Adder m_639 ( // @[MUL.scala 124:19]
    .io_in_0(m_639_io_in_0),
    .io_in_1(m_639_io_in_1),
    .io_out_0(m_639_io_out_0),
    .io_out_1(m_639_io_out_1)
  );
  Half_Adder m_640 ( // @[MUL.scala 124:19]
    .io_in_0(m_640_io_in_0),
    .io_in_1(m_640_io_in_1),
    .io_out_0(m_640_io_out_0),
    .io_out_1(m_640_io_out_1)
  );
  Half_Adder m_641 ( // @[MUL.scala 124:19]
    .io_in_0(m_641_io_in_0),
    .io_in_1(m_641_io_in_1),
    .io_out_0(m_641_io_out_0),
    .io_out_1(m_641_io_out_1)
  );
  Half_Adder m_642 ( // @[MUL.scala 124:19]
    .io_in_0(m_642_io_in_0),
    .io_in_1(m_642_io_in_1),
    .io_out_0(m_642_io_out_0),
    .io_out_1(m_642_io_out_1)
  );
  Half_Adder m_643 ( // @[MUL.scala 124:19]
    .io_in_0(m_643_io_in_0),
    .io_in_1(m_643_io_in_1),
    .io_out_0(m_643_io_out_0),
    .io_out_1(m_643_io_out_1)
  );
  Half_Adder m_644 ( // @[MUL.scala 124:19]
    .io_in_0(m_644_io_in_0),
    .io_in_1(m_644_io_in_1),
    .io_out_0(m_644_io_out_0),
    .io_out_1(m_644_io_out_1)
  );
  Half_Adder m_645 ( // @[MUL.scala 124:19]
    .io_in_0(m_645_io_in_0),
    .io_in_1(m_645_io_in_1),
    .io_out_0(m_645_io_out_0),
    .io_out_1(m_645_io_out_1)
  );
  Half_Adder m_646 ( // @[MUL.scala 124:19]
    .io_in_0(m_646_io_in_0),
    .io_in_1(m_646_io_in_1),
    .io_out_0(m_646_io_out_0),
    .io_out_1(m_646_io_out_1)
  );
  Half_Adder m_647 ( // @[MUL.scala 124:19]
    .io_in_0(m_647_io_in_0),
    .io_in_1(m_647_io_in_1),
    .io_out_0(m_647_io_out_0),
    .io_out_1(m_647_io_out_1)
  );
  Half_Adder m_648 ( // @[MUL.scala 124:19]
    .io_in_0(m_648_io_in_0),
    .io_in_1(m_648_io_in_1),
    .io_out_0(m_648_io_out_0),
    .io_out_1(m_648_io_out_1)
  );
  Half_Adder m_649 ( // @[MUL.scala 124:19]
    .io_in_0(m_649_io_in_0),
    .io_in_1(m_649_io_in_1),
    .io_out_0(m_649_io_out_0),
    .io_out_1(m_649_io_out_1)
  );
  Half_Adder m_650 ( // @[MUL.scala 124:19]
    .io_in_0(m_650_io_in_0),
    .io_in_1(m_650_io_in_1),
    .io_out_0(m_650_io_out_0),
    .io_out_1(m_650_io_out_1)
  );
  Half_Adder m_651 ( // @[MUL.scala 124:19]
    .io_in_0(m_651_io_in_0),
    .io_in_1(m_651_io_in_1),
    .io_out_0(m_651_io_out_0),
    .io_out_1(m_651_io_out_1)
  );
  Half_Adder m_652 ( // @[MUL.scala 124:19]
    .io_in_0(m_652_io_in_0),
    .io_in_1(m_652_io_in_1),
    .io_out_0(m_652_io_out_0),
    .io_out_1(m_652_io_out_1)
  );
  Half_Adder m_653 ( // @[MUL.scala 124:19]
    .io_in_0(m_653_io_in_0),
    .io_in_1(m_653_io_in_1),
    .io_out_0(m_653_io_out_0),
    .io_out_1(m_653_io_out_1)
  );
  Half_Adder m_654 ( // @[MUL.scala 124:19]
    .io_in_0(m_654_io_in_0),
    .io_in_1(m_654_io_in_1),
    .io_out_0(m_654_io_out_0),
    .io_out_1(m_654_io_out_1)
  );
  Half_Adder m_655 ( // @[MUL.scala 124:19]
    .io_in_0(m_655_io_in_0),
    .io_in_1(m_655_io_in_1),
    .io_out_0(m_655_io_out_0),
    .io_out_1(m_655_io_out_1)
  );
  Half_Adder m_656 ( // @[MUL.scala 124:19]
    .io_in_0(m_656_io_in_0),
    .io_in_1(m_656_io_in_1),
    .io_out_0(m_656_io_out_0),
    .io_out_1(m_656_io_out_1)
  );
  Half_Adder m_657 ( // @[MUL.scala 124:19]
    .io_in_0(m_657_io_in_0),
    .io_in_1(m_657_io_in_1),
    .io_out_0(m_657_io_out_0),
    .io_out_1(m_657_io_out_1)
  );
  Half_Adder m_658 ( // @[MUL.scala 124:19]
    .io_in_0(m_658_io_in_0),
    .io_in_1(m_658_io_in_1),
    .io_out_0(m_658_io_out_0),
    .io_out_1(m_658_io_out_1)
  );
  Half_Adder m_659 ( // @[MUL.scala 124:19]
    .io_in_0(m_659_io_in_0),
    .io_in_1(m_659_io_in_1),
    .io_out_0(m_659_io_out_0),
    .io_out_1(m_659_io_out_1)
  );
  Half_Adder m_660 ( // @[MUL.scala 124:19]
    .io_in_0(m_660_io_in_0),
    .io_in_1(m_660_io_in_1),
    .io_out_0(m_660_io_out_0),
    .io_out_1(m_660_io_out_1)
  );
  Adder m_661 ( // @[MUL.scala 102:19]
    .io_x1(m_661_io_x1),
    .io_x2(m_661_io_x2),
    .io_x3(m_661_io_x3),
    .io_s(m_661_io_s),
    .io_cout(m_661_io_cout)
  );
  Adder m_662 ( // @[MUL.scala 102:19]
    .io_x1(m_662_io_x1),
    .io_x2(m_662_io_x2),
    .io_x3(m_662_io_x3),
    .io_s(m_662_io_s),
    .io_cout(m_662_io_cout)
  );
  Adder m_663 ( // @[MUL.scala 102:19]
    .io_x1(m_663_io_x1),
    .io_x2(m_663_io_x2),
    .io_x3(m_663_io_x3),
    .io_s(m_663_io_s),
    .io_cout(m_663_io_cout)
  );
  Adder m_664 ( // @[MUL.scala 102:19]
    .io_x1(m_664_io_x1),
    .io_x2(m_664_io_x2),
    .io_x3(m_664_io_x3),
    .io_s(m_664_io_s),
    .io_cout(m_664_io_cout)
  );
  Adder m_665 ( // @[MUL.scala 102:19]
    .io_x1(m_665_io_x1),
    .io_x2(m_665_io_x2),
    .io_x3(m_665_io_x3),
    .io_s(m_665_io_s),
    .io_cout(m_665_io_cout)
  );
  Adder m_666 ( // @[MUL.scala 102:19]
    .io_x1(m_666_io_x1),
    .io_x2(m_666_io_x2),
    .io_x3(m_666_io_x3),
    .io_s(m_666_io_s),
    .io_cout(m_666_io_cout)
  );
  Adder m_667 ( // @[MUL.scala 102:19]
    .io_x1(m_667_io_x1),
    .io_x2(m_667_io_x2),
    .io_x3(m_667_io_x3),
    .io_s(m_667_io_s),
    .io_cout(m_667_io_cout)
  );
  Adder m_668 ( // @[MUL.scala 102:19]
    .io_x1(m_668_io_x1),
    .io_x2(m_668_io_x2),
    .io_x3(m_668_io_x3),
    .io_s(m_668_io_s),
    .io_cout(m_668_io_cout)
  );
  Adder m_669 ( // @[MUL.scala 102:19]
    .io_x1(m_669_io_x1),
    .io_x2(m_669_io_x2),
    .io_x3(m_669_io_x3),
    .io_s(m_669_io_s),
    .io_cout(m_669_io_cout)
  );
  Adder m_670 ( // @[MUL.scala 102:19]
    .io_x1(m_670_io_x1),
    .io_x2(m_670_io_x2),
    .io_x3(m_670_io_x3),
    .io_s(m_670_io_s),
    .io_cout(m_670_io_cout)
  );
  Adder m_671 ( // @[MUL.scala 102:19]
    .io_x1(m_671_io_x1),
    .io_x2(m_671_io_x2),
    .io_x3(m_671_io_x3),
    .io_s(m_671_io_s),
    .io_cout(m_671_io_cout)
  );
  Adder m_672 ( // @[MUL.scala 102:19]
    .io_x1(m_672_io_x1),
    .io_x2(m_672_io_x2),
    .io_x3(m_672_io_x3),
    .io_s(m_672_io_s),
    .io_cout(m_672_io_cout)
  );
  Adder m_673 ( // @[MUL.scala 102:19]
    .io_x1(m_673_io_x1),
    .io_x2(m_673_io_x2),
    .io_x3(m_673_io_x3),
    .io_s(m_673_io_s),
    .io_cout(m_673_io_cout)
  );
  Adder m_674 ( // @[MUL.scala 102:19]
    .io_x1(m_674_io_x1),
    .io_x2(m_674_io_x2),
    .io_x3(m_674_io_x3),
    .io_s(m_674_io_s),
    .io_cout(m_674_io_cout)
  );
  Adder m_675 ( // @[MUL.scala 102:19]
    .io_x1(m_675_io_x1),
    .io_x2(m_675_io_x2),
    .io_x3(m_675_io_x3),
    .io_s(m_675_io_s),
    .io_cout(m_675_io_cout)
  );
  Adder m_676 ( // @[MUL.scala 102:19]
    .io_x1(m_676_io_x1),
    .io_x2(m_676_io_x2),
    .io_x3(m_676_io_x3),
    .io_s(m_676_io_s),
    .io_cout(m_676_io_cout)
  );
  Adder m_677 ( // @[MUL.scala 102:19]
    .io_x1(m_677_io_x1),
    .io_x2(m_677_io_x2),
    .io_x3(m_677_io_x3),
    .io_s(m_677_io_s),
    .io_cout(m_677_io_cout)
  );
  Adder m_678 ( // @[MUL.scala 102:19]
    .io_x1(m_678_io_x1),
    .io_x2(m_678_io_x2),
    .io_x3(m_678_io_x3),
    .io_s(m_678_io_s),
    .io_cout(m_678_io_cout)
  );
  Half_Adder m_679 ( // @[MUL.scala 124:19]
    .io_in_0(m_679_io_in_0),
    .io_in_1(m_679_io_in_1),
    .io_out_0(m_679_io_out_0),
    .io_out_1(m_679_io_out_1)
  );
  Half_Adder m_680 ( // @[MUL.scala 124:19]
    .io_in_0(m_680_io_in_0),
    .io_in_1(m_680_io_in_1),
    .io_out_0(m_680_io_out_0),
    .io_out_1(m_680_io_out_1)
  );
  Half_Adder m_681 ( // @[MUL.scala 124:19]
    .io_in_0(m_681_io_in_0),
    .io_in_1(m_681_io_in_1),
    .io_out_0(m_681_io_out_0),
    .io_out_1(m_681_io_out_1)
  );
  Half_Adder m_682 ( // @[MUL.scala 124:19]
    .io_in_0(m_682_io_in_0),
    .io_in_1(m_682_io_in_1),
    .io_out_0(m_682_io_out_0),
    .io_out_1(m_682_io_out_1)
  );
  Half_Adder m_683 ( // @[MUL.scala 124:19]
    .io_in_0(m_683_io_in_0),
    .io_in_1(m_683_io_in_1),
    .io_out_0(m_683_io_out_0),
    .io_out_1(m_683_io_out_1)
  );
  Half_Adder m_684 ( // @[MUL.scala 124:19]
    .io_in_0(m_684_io_in_0),
    .io_in_1(m_684_io_in_1),
    .io_out_0(m_684_io_out_0),
    .io_out_1(m_684_io_out_1)
  );
  Half_Adder m_685 ( // @[MUL.scala 124:19]
    .io_in_0(m_685_io_in_0),
    .io_in_1(m_685_io_in_1),
    .io_out_0(m_685_io_out_0),
    .io_out_1(m_685_io_out_1)
  );
  Half_Adder m_686 ( // @[MUL.scala 124:19]
    .io_in_0(m_686_io_in_0),
    .io_in_1(m_686_io_in_1),
    .io_out_0(m_686_io_out_0),
    .io_out_1(m_686_io_out_1)
  );
  Half_Adder m_687 ( // @[MUL.scala 124:19]
    .io_in_0(m_687_io_in_0),
    .io_in_1(m_687_io_in_1),
    .io_out_0(m_687_io_out_0),
    .io_out_1(m_687_io_out_1)
  );
  Half_Adder m_688 ( // @[MUL.scala 124:19]
    .io_in_0(m_688_io_in_0),
    .io_in_1(m_688_io_in_1),
    .io_out_0(m_688_io_out_0),
    .io_out_1(m_688_io_out_1)
  );
  Half_Adder m_689 ( // @[MUL.scala 124:19]
    .io_in_0(m_689_io_in_0),
    .io_in_1(m_689_io_in_1),
    .io_out_0(m_689_io_out_0),
    .io_out_1(m_689_io_out_1)
  );
  Half_Adder m_690 ( // @[MUL.scala 124:19]
    .io_in_0(m_690_io_in_0),
    .io_in_1(m_690_io_in_1),
    .io_out_0(m_690_io_out_0),
    .io_out_1(m_690_io_out_1)
  );
  Half_Adder m_691 ( // @[MUL.scala 124:19]
    .io_in_0(m_691_io_in_0),
    .io_in_1(m_691_io_in_1),
    .io_out_0(m_691_io_out_0),
    .io_out_1(m_691_io_out_1)
  );
  Half_Adder m_692 ( // @[MUL.scala 124:19]
    .io_in_0(m_692_io_in_0),
    .io_in_1(m_692_io_in_1),
    .io_out_0(m_692_io_out_0),
    .io_out_1(m_692_io_out_1)
  );
  Half_Adder m_693 ( // @[MUL.scala 124:19]
    .io_in_0(m_693_io_in_0),
    .io_in_1(m_693_io_in_1),
    .io_out_0(m_693_io_out_0),
    .io_out_1(m_693_io_out_1)
  );
  Half_Adder m_694 ( // @[MUL.scala 124:19]
    .io_in_0(m_694_io_in_0),
    .io_in_1(m_694_io_in_1),
    .io_out_0(m_694_io_out_0),
    .io_out_1(m_694_io_out_1)
  );
  Half_Adder m_695 ( // @[MUL.scala 124:19]
    .io_in_0(m_695_io_in_0),
    .io_in_1(m_695_io_in_1),
    .io_out_0(m_695_io_out_0),
    .io_out_1(m_695_io_out_1)
  );
  Half_Adder m_696 ( // @[MUL.scala 124:19]
    .io_in_0(m_696_io_in_0),
    .io_in_1(m_696_io_in_1),
    .io_out_0(m_696_io_out_0),
    .io_out_1(m_696_io_out_1)
  );
  Half_Adder m_697 ( // @[MUL.scala 124:19]
    .io_in_0(m_697_io_in_0),
    .io_in_1(m_697_io_in_1),
    .io_out_0(m_697_io_out_0),
    .io_out_1(m_697_io_out_1)
  );
  Half_Adder m_698 ( // @[MUL.scala 124:19]
    .io_in_0(m_698_io_in_0),
    .io_in_1(m_698_io_in_1),
    .io_out_0(m_698_io_out_0),
    .io_out_1(m_698_io_out_1)
  );
  Half_Adder m_699 ( // @[MUL.scala 124:19]
    .io_in_0(m_699_io_in_0),
    .io_in_1(m_699_io_in_1),
    .io_out_0(m_699_io_out_0),
    .io_out_1(m_699_io_out_1)
  );
  Half_Adder m_700 ( // @[MUL.scala 124:19]
    .io_in_0(m_700_io_in_0),
    .io_in_1(m_700_io_in_1),
    .io_out_0(m_700_io_out_0),
    .io_out_1(m_700_io_out_1)
  );
  Half_Adder m_701 ( // @[MUL.scala 124:19]
    .io_in_0(m_701_io_in_0),
    .io_in_1(m_701_io_in_1),
    .io_out_0(m_701_io_out_0),
    .io_out_1(m_701_io_out_1)
  );
  assign io_in_ready = 1'h1; // @[MUL.scala 356:15]
  assign io_out_valid = count == 8'h2; // @[MUL.scala 345:17]
  assign io_out_bits_result_result_hi = result[63:32]; // @[MUL.scala 353:41]
  assign io_out_bits_result_result_lo = result[31:0]; // @[MUL.scala 354:40]
  assign m_io_y_3 = src1[2:0]; // @[MUL.scala 313:56]
  assign m_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_1_io_y_3 = src1[4:2]; // @[MUL.scala 313:56]
  assign m_1_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_2_io_y_3 = src1[6:4]; // @[MUL.scala 313:56]
  assign m_2_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_3_io_y_3 = src1[8:6]; // @[MUL.scala 313:56]
  assign m_3_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_4_io_y_3 = src1[10:8]; // @[MUL.scala 313:56]
  assign m_4_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_5_io_y_3 = src1[12:10]; // @[MUL.scala 313:56]
  assign m_5_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_6_io_y_3 = src1[14:12]; // @[MUL.scala 313:56]
  assign m_6_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_7_io_y_3 = src1[16:14]; // @[MUL.scala 313:56]
  assign m_7_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_8_io_y_3 = src1[18:16]; // @[MUL.scala 313:56]
  assign m_8_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_9_io_y_3 = src1[20:18]; // @[MUL.scala 313:56]
  assign m_9_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_10_io_y_3 = src1[22:20]; // @[MUL.scala 313:56]
  assign m_10_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_11_io_y_3 = src1[24:22]; // @[MUL.scala 313:56]
  assign m_11_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_12_io_y_3 = src1[26:24]; // @[MUL.scala 313:56]
  assign m_12_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_13_io_y_3 = src1[28:26]; // @[MUL.scala 313:56]
  assign m_13_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_14_io_y_3 = src1[30:28]; // @[MUL.scala 313:56]
  assign m_14_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_15_io_y_3 = src1[32:30]; // @[MUL.scala 313:56]
  assign m_15_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_16_io_y_3 = src1[34:32]; // @[MUL.scala 313:56]
  assign m_16_io_x = _src2_T_6 | _src2_T_5; // @[Mux.scala 27:73]
  assign m_17_io_in_0 = r; // @[MUL.scala 125:16]
  assign m_17_io_in_1 = r_1; // @[MUL.scala 126:16]
  assign m_18_io_in_0 = r_2; // @[MUL.scala 125:16]
  assign m_18_io_in_1 = r_3; // @[MUL.scala 126:16]
  assign m_19_io_x1 = r_4; // @[MUL.scala 103:13]
  assign m_19_io_x2 = r_5; // @[MUL.scala 104:13]
  assign m_19_io_x3 = r_6; // @[MUL.scala 105:13]
  assign m_20_io_x1 = r_7; // @[MUL.scala 103:13]
  assign m_20_io_x2 = r_8; // @[MUL.scala 104:13]
  assign m_20_io_x3 = r_9; // @[MUL.scala 105:13]
  assign m_21_io_x1 = r_10; // @[MUL.scala 103:13]
  assign m_21_io_x2 = r_11; // @[MUL.scala 104:13]
  assign m_21_io_x3 = r_12; // @[MUL.scala 105:13]
  assign m_22_io_x1 = r_14; // @[MUL.scala 103:13]
  assign m_22_io_x2 = r_15; // @[MUL.scala 104:13]
  assign m_22_io_x3 = r_16; // @[MUL.scala 105:13]
  assign m_23_io_x1 = r_18; // @[MUL.scala 103:13]
  assign m_23_io_x2 = r_19; // @[MUL.scala 104:13]
  assign m_23_io_x3 = r_20; // @[MUL.scala 105:13]
  assign m_24_io_in_0 = r_21; // @[MUL.scala 125:16]
  assign m_24_io_in_1 = r_22; // @[MUL.scala 126:16]
  assign m_25_io_x1 = r_23; // @[MUL.scala 103:13]
  assign m_25_io_x2 = r_24; // @[MUL.scala 104:13]
  assign m_25_io_x3 = r_25; // @[MUL.scala 105:13]
  assign m_26_io_in_0 = r_26; // @[MUL.scala 125:16]
  assign m_26_io_in_1 = r_27; // @[MUL.scala 126:16]
  assign m_27_io_x1 = r_28; // @[MUL.scala 103:13]
  assign m_27_io_x2 = r_29; // @[MUL.scala 104:13]
  assign m_27_io_x3 = r_30; // @[MUL.scala 105:13]
  assign m_28_io_x1 = r_31; // @[MUL.scala 103:13]
  assign m_28_io_x2 = r_32; // @[MUL.scala 104:13]
  assign m_28_io_x3 = r_33; // @[MUL.scala 105:13]
  assign m_29_io_x1 = r_34; // @[MUL.scala 103:13]
  assign m_29_io_x2 = r_35; // @[MUL.scala 104:13]
  assign m_29_io_x3 = r_36; // @[MUL.scala 105:13]
  assign m_30_io_x1 = r_37; // @[MUL.scala 103:13]
  assign m_30_io_x2 = r_38; // @[MUL.scala 104:13]
  assign m_30_io_x3 = r_39; // @[MUL.scala 105:13]
  assign m_31_io_x1 = r_40; // @[MUL.scala 103:13]
  assign m_31_io_x2 = r_41; // @[MUL.scala 104:13]
  assign m_31_io_x3 = r_42; // @[MUL.scala 105:13]
  assign m_32_io_x1 = r_43; // @[MUL.scala 103:13]
  assign m_32_io_x2 = r_44; // @[MUL.scala 104:13]
  assign m_32_io_x3 = r_45; // @[MUL.scala 105:13]
  assign m_33_io_x1 = r_47; // @[MUL.scala 103:13]
  assign m_33_io_x2 = r_48; // @[MUL.scala 104:13]
  assign m_33_io_x3 = r_49; // @[MUL.scala 105:13]
  assign m_34_io_x1 = r_50; // @[MUL.scala 103:13]
  assign m_34_io_x2 = r_51; // @[MUL.scala 104:13]
  assign m_34_io_x3 = r_52; // @[MUL.scala 105:13]
  assign m_35_io_x1 = r_54; // @[MUL.scala 103:13]
  assign m_35_io_x2 = r_55; // @[MUL.scala 104:13]
  assign m_35_io_x3 = r_56; // @[MUL.scala 105:13]
  assign m_36_io_x1 = r_57; // @[MUL.scala 103:13]
  assign m_36_io_x2 = r_58; // @[MUL.scala 104:13]
  assign m_36_io_x3 = r_59; // @[MUL.scala 105:13]
  assign m_37_io_in_0 = r_60; // @[MUL.scala 125:16]
  assign m_37_io_in_1 = r_61; // @[MUL.scala 126:16]
  assign m_38_io_x1 = r_62; // @[MUL.scala 103:13]
  assign m_38_io_x2 = r_63; // @[MUL.scala 104:13]
  assign m_38_io_x3 = r_64; // @[MUL.scala 105:13]
  assign m_39_io_x1 = r_65; // @[MUL.scala 103:13]
  assign m_39_io_x2 = r_66; // @[MUL.scala 104:13]
  assign m_39_io_x3 = r_67; // @[MUL.scala 105:13]
  assign m_40_io_in_0 = r_68; // @[MUL.scala 125:16]
  assign m_40_io_in_1 = r_69; // @[MUL.scala 126:16]
  assign m_41_io_x1 = r_70; // @[MUL.scala 103:13]
  assign m_41_io_x2 = r_71; // @[MUL.scala 104:13]
  assign m_41_io_x3 = r_72; // @[MUL.scala 105:13]
  assign m_42_io_x1 = r_73; // @[MUL.scala 103:13]
  assign m_42_io_x2 = r_74; // @[MUL.scala 104:13]
  assign m_42_io_x3 = r_75; // @[MUL.scala 105:13]
  assign m_43_io_x1 = r_76; // @[MUL.scala 103:13]
  assign m_43_io_x2 = r_77; // @[MUL.scala 104:13]
  assign m_43_io_x3 = r_78; // @[MUL.scala 105:13]
  assign m_44_io_x1 = r_79; // @[MUL.scala 103:13]
  assign m_44_io_x2 = r_80; // @[MUL.scala 104:13]
  assign m_44_io_x3 = r_81; // @[MUL.scala 105:13]
  assign m_45_io_x1 = r_82; // @[MUL.scala 103:13]
  assign m_45_io_x2 = r_83; // @[MUL.scala 104:13]
  assign m_45_io_x3 = r_84; // @[MUL.scala 105:13]
  assign m_46_io_x1 = r_85; // @[MUL.scala 103:13]
  assign m_46_io_x2 = r_86; // @[MUL.scala 104:13]
  assign m_46_io_x3 = r_87; // @[MUL.scala 105:13]
  assign m_47_io_x1 = r_88; // @[MUL.scala 103:13]
  assign m_47_io_x2 = r_89; // @[MUL.scala 104:13]
  assign m_47_io_x3 = r_90; // @[MUL.scala 105:13]
  assign m_48_io_x1 = r_91; // @[MUL.scala 103:13]
  assign m_48_io_x2 = r_92; // @[MUL.scala 104:13]
  assign m_48_io_x3 = r_93; // @[MUL.scala 105:13]
  assign m_49_io_x1 = r_94; // @[MUL.scala 103:13]
  assign m_49_io_x2 = r_95; // @[MUL.scala 104:13]
  assign m_49_io_x3 = r_96; // @[MUL.scala 105:13]
  assign m_50_io_x1 = r_98; // @[MUL.scala 103:13]
  assign m_50_io_x2 = r_99; // @[MUL.scala 104:13]
  assign m_50_io_x3 = r_100; // @[MUL.scala 105:13]
  assign m_51_io_x1 = r_101; // @[MUL.scala 103:13]
  assign m_51_io_x2 = r_102; // @[MUL.scala 104:13]
  assign m_51_io_x3 = r_103; // @[MUL.scala 105:13]
  assign m_52_io_x1 = r_104; // @[MUL.scala 103:13]
  assign m_52_io_x2 = r_105; // @[MUL.scala 104:13]
  assign m_52_io_x3 = r_106; // @[MUL.scala 105:13]
  assign m_53_io_x1 = r_108; // @[MUL.scala 103:13]
  assign m_53_io_x2 = r_109; // @[MUL.scala 104:13]
  assign m_53_io_x3 = r_110; // @[MUL.scala 105:13]
  assign m_54_io_x1 = r_111; // @[MUL.scala 103:13]
  assign m_54_io_x2 = r_112; // @[MUL.scala 104:13]
  assign m_54_io_x3 = r_113; // @[MUL.scala 105:13]
  assign m_55_io_x1 = r_114; // @[MUL.scala 103:13]
  assign m_55_io_x2 = r_115; // @[MUL.scala 104:13]
  assign m_55_io_x3 = r_116; // @[MUL.scala 105:13]
  assign m_56_io_in_0 = r_117; // @[MUL.scala 125:16]
  assign m_56_io_in_1 = r_118; // @[MUL.scala 126:16]
  assign m_57_io_x1 = r_119; // @[MUL.scala 103:13]
  assign m_57_io_x2 = r_120; // @[MUL.scala 104:13]
  assign m_57_io_x3 = r_121; // @[MUL.scala 105:13]
  assign m_58_io_x1 = r_122; // @[MUL.scala 103:13]
  assign m_58_io_x2 = r_123; // @[MUL.scala 104:13]
  assign m_58_io_x3 = r_124; // @[MUL.scala 105:13]
  assign m_59_io_x1 = r_125; // @[MUL.scala 103:13]
  assign m_59_io_x2 = r_126; // @[MUL.scala 104:13]
  assign m_59_io_x3 = r_127; // @[MUL.scala 105:13]
  assign m_60_io_in_0 = r_128; // @[MUL.scala 125:16]
  assign m_60_io_in_1 = r_129; // @[MUL.scala 126:16]
  assign m_61_io_x1 = r_130; // @[MUL.scala 103:13]
  assign m_61_io_x2 = r_131; // @[MUL.scala 104:13]
  assign m_61_io_x3 = r_132; // @[MUL.scala 105:13]
  assign m_62_io_x1 = r_133; // @[MUL.scala 103:13]
  assign m_62_io_x2 = r_134; // @[MUL.scala 104:13]
  assign m_62_io_x3 = r_135; // @[MUL.scala 105:13]
  assign m_63_io_x1 = r_136; // @[MUL.scala 103:13]
  assign m_63_io_x2 = r_137; // @[MUL.scala 104:13]
  assign m_63_io_x3 = r_138; // @[MUL.scala 105:13]
  assign m_64_io_x1 = r_139; // @[MUL.scala 103:13]
  assign m_64_io_x2 = r_140; // @[MUL.scala 104:13]
  assign m_64_io_x3 = r_141; // @[MUL.scala 105:13]
  assign m_65_io_x1 = r_142; // @[MUL.scala 103:13]
  assign m_65_io_x2 = r_143; // @[MUL.scala 104:13]
  assign m_65_io_x3 = r_144; // @[MUL.scala 105:13]
  assign m_66_io_x1 = r_145; // @[MUL.scala 103:13]
  assign m_66_io_x2 = r_146; // @[MUL.scala 104:13]
  assign m_66_io_x3 = r_147; // @[MUL.scala 105:13]
  assign m_67_io_x1 = r_148; // @[MUL.scala 103:13]
  assign m_67_io_x2 = r_149; // @[MUL.scala 104:13]
  assign m_67_io_x3 = r_150; // @[MUL.scala 105:13]
  assign m_68_io_x1 = r_151; // @[MUL.scala 103:13]
  assign m_68_io_x2 = r_152; // @[MUL.scala 104:13]
  assign m_68_io_x3 = r_153; // @[MUL.scala 105:13]
  assign m_69_io_x1 = r_154; // @[MUL.scala 103:13]
  assign m_69_io_x2 = r_155; // @[MUL.scala 104:13]
  assign m_69_io_x3 = r_156; // @[MUL.scala 105:13]
  assign m_70_io_x1 = r_157; // @[MUL.scala 103:13]
  assign m_70_io_x2 = r_158; // @[MUL.scala 104:13]
  assign m_70_io_x3 = r_159; // @[MUL.scala 105:13]
  assign m_71_io_x1 = r_160; // @[MUL.scala 103:13]
  assign m_71_io_x2 = r_161; // @[MUL.scala 104:13]
  assign m_71_io_x3 = r_162; // @[MUL.scala 105:13]
  assign m_72_io_x1 = r_163; // @[MUL.scala 103:13]
  assign m_72_io_x2 = r_164; // @[MUL.scala 104:13]
  assign m_72_io_x3 = r_165; // @[MUL.scala 105:13]
  assign m_73_io_x1 = r_167; // @[MUL.scala 103:13]
  assign m_73_io_x2 = r_168; // @[MUL.scala 104:13]
  assign m_73_io_x3 = r_169; // @[MUL.scala 105:13]
  assign m_74_io_x1 = r_170; // @[MUL.scala 103:13]
  assign m_74_io_x2 = r_171; // @[MUL.scala 104:13]
  assign m_74_io_x3 = r_172; // @[MUL.scala 105:13]
  assign m_75_io_x1 = r_173; // @[MUL.scala 103:13]
  assign m_75_io_x2 = r_174; // @[MUL.scala 104:13]
  assign m_75_io_x3 = r_175; // @[MUL.scala 105:13]
  assign m_76_io_x1 = r_176; // @[MUL.scala 103:13]
  assign m_76_io_x2 = r_177; // @[MUL.scala 104:13]
  assign m_76_io_x3 = r_178; // @[MUL.scala 105:13]
  assign m_77_io_x1 = r_180; // @[MUL.scala 103:13]
  assign m_77_io_x2 = r_181; // @[MUL.scala 104:13]
  assign m_77_io_x3 = r_182; // @[MUL.scala 105:13]
  assign m_78_io_x1 = r_183; // @[MUL.scala 103:13]
  assign m_78_io_x2 = r_184; // @[MUL.scala 104:13]
  assign m_78_io_x3 = r_185; // @[MUL.scala 105:13]
  assign m_79_io_x1 = r_186; // @[MUL.scala 103:13]
  assign m_79_io_x2 = r_187; // @[MUL.scala 104:13]
  assign m_79_io_x3 = r_188; // @[MUL.scala 105:13]
  assign m_80_io_x1 = r_189; // @[MUL.scala 103:13]
  assign m_80_io_x2 = r_190; // @[MUL.scala 104:13]
  assign m_80_io_x3 = r_191; // @[MUL.scala 105:13]
  assign m_81_io_in_0 = r_192; // @[MUL.scala 125:16]
  assign m_81_io_in_1 = r_193; // @[MUL.scala 126:16]
  assign m_82_io_x1 = r_194; // @[MUL.scala 103:13]
  assign m_82_io_x2 = r_195; // @[MUL.scala 104:13]
  assign m_82_io_x3 = r_196; // @[MUL.scala 105:13]
  assign m_83_io_x1 = r_197; // @[MUL.scala 103:13]
  assign m_83_io_x2 = r_198; // @[MUL.scala 104:13]
  assign m_83_io_x3 = r_199; // @[MUL.scala 105:13]
  assign m_84_io_x1 = r_200; // @[MUL.scala 103:13]
  assign m_84_io_x2 = r_201; // @[MUL.scala 104:13]
  assign m_84_io_x3 = r_202; // @[MUL.scala 105:13]
  assign m_85_io_x1 = r_203; // @[MUL.scala 103:13]
  assign m_85_io_x2 = r_204; // @[MUL.scala 104:13]
  assign m_85_io_x3 = r_205; // @[MUL.scala 105:13]
  assign m_86_io_in_0 = r_206; // @[MUL.scala 125:16]
  assign m_86_io_in_1 = r_207; // @[MUL.scala 126:16]
  assign m_87_io_x1 = r_208; // @[MUL.scala 103:13]
  assign m_87_io_x2 = r_209; // @[MUL.scala 104:13]
  assign m_87_io_x3 = r_210; // @[MUL.scala 105:13]
  assign m_88_io_x1 = r_211; // @[MUL.scala 103:13]
  assign m_88_io_x2 = r_212; // @[MUL.scala 104:13]
  assign m_88_io_x3 = r_213; // @[MUL.scala 105:13]
  assign m_89_io_x1 = r_214; // @[MUL.scala 103:13]
  assign m_89_io_x2 = r_215; // @[MUL.scala 104:13]
  assign m_89_io_x3 = r_216; // @[MUL.scala 105:13]
  assign m_90_io_x1 = r_217; // @[MUL.scala 103:13]
  assign m_90_io_x2 = r_218; // @[MUL.scala 104:13]
  assign m_90_io_x3 = r_219; // @[MUL.scala 105:13]
  assign m_91_io_x1 = r_220; // @[MUL.scala 103:13]
  assign m_91_io_x2 = r_221; // @[MUL.scala 104:13]
  assign m_91_io_x3 = r_222; // @[MUL.scala 105:13]
  assign m_92_io_x1 = r_223; // @[MUL.scala 103:13]
  assign m_92_io_x2 = r_224; // @[MUL.scala 104:13]
  assign m_92_io_x3 = r_225; // @[MUL.scala 105:13]
  assign m_93_io_x1 = r_226; // @[MUL.scala 103:13]
  assign m_93_io_x2 = r_227; // @[MUL.scala 104:13]
  assign m_93_io_x3 = r_228; // @[MUL.scala 105:13]
  assign m_94_io_x1 = r_229; // @[MUL.scala 103:13]
  assign m_94_io_x2 = r_230; // @[MUL.scala 104:13]
  assign m_94_io_x3 = r_231; // @[MUL.scala 105:13]
  assign m_95_io_x1 = r_232; // @[MUL.scala 103:13]
  assign m_95_io_x2 = r_233; // @[MUL.scala 104:13]
  assign m_95_io_x3 = r_234; // @[MUL.scala 105:13]
  assign m_96_io_x1 = r_235; // @[MUL.scala 103:13]
  assign m_96_io_x2 = r_236; // @[MUL.scala 104:13]
  assign m_96_io_x3 = r_237; // @[MUL.scala 105:13]
  assign m_97_io_x1 = r_238; // @[MUL.scala 103:13]
  assign m_97_io_x2 = r_239; // @[MUL.scala 104:13]
  assign m_97_io_x3 = r_240; // @[MUL.scala 105:13]
  assign m_98_io_x1 = r_241; // @[MUL.scala 103:13]
  assign m_98_io_x2 = r_242; // @[MUL.scala 104:13]
  assign m_98_io_x3 = r_243; // @[MUL.scala 105:13]
  assign m_99_io_x1 = r_244; // @[MUL.scala 103:13]
  assign m_99_io_x2 = r_245; // @[MUL.scala 104:13]
  assign m_99_io_x3 = r_246; // @[MUL.scala 105:13]
  assign m_100_io_x1 = r_247; // @[MUL.scala 103:13]
  assign m_100_io_x2 = r_248; // @[MUL.scala 104:13]
  assign m_100_io_x3 = r_249; // @[MUL.scala 105:13]
  assign m_101_io_x1 = r_250; // @[MUL.scala 103:13]
  assign m_101_io_x2 = r_251; // @[MUL.scala 104:13]
  assign m_101_io_x3 = r_252; // @[MUL.scala 105:13]
  assign m_102_io_x1 = r_254; // @[MUL.scala 103:13]
  assign m_102_io_x2 = r_255; // @[MUL.scala 104:13]
  assign m_102_io_x3 = r_256; // @[MUL.scala 105:13]
  assign m_103_io_x1 = r_257; // @[MUL.scala 103:13]
  assign m_103_io_x2 = r_258; // @[MUL.scala 104:13]
  assign m_103_io_x3 = r_259; // @[MUL.scala 105:13]
  assign m_104_io_x1 = r_260; // @[MUL.scala 103:13]
  assign m_104_io_x2 = r_261; // @[MUL.scala 104:13]
  assign m_104_io_x3 = r_262; // @[MUL.scala 105:13]
  assign m_105_io_x1 = r_263; // @[MUL.scala 103:13]
  assign m_105_io_x2 = r_264; // @[MUL.scala 104:13]
  assign m_105_io_x3 = r_265; // @[MUL.scala 105:13]
  assign m_106_io_x1 = r_266; // @[MUL.scala 103:13]
  assign m_106_io_x2 = r_267; // @[MUL.scala 104:13]
  assign m_106_io_x3 = r_268; // @[MUL.scala 105:13]
  assign m_107_io_x1 = r_270; // @[MUL.scala 103:13]
  assign m_107_io_x2 = r_271; // @[MUL.scala 104:13]
  assign m_107_io_x3 = r_272; // @[MUL.scala 105:13]
  assign m_108_io_x1 = r_273; // @[MUL.scala 103:13]
  assign m_108_io_x2 = r_274; // @[MUL.scala 104:13]
  assign m_108_io_x3 = r_275; // @[MUL.scala 105:13]
  assign m_109_io_x1 = r_276; // @[MUL.scala 103:13]
  assign m_109_io_x2 = r_277; // @[MUL.scala 104:13]
  assign m_109_io_x3 = r_278; // @[MUL.scala 105:13]
  assign m_110_io_x1 = r_279; // @[MUL.scala 103:13]
  assign m_110_io_x2 = r_280; // @[MUL.scala 104:13]
  assign m_110_io_x3 = r_281; // @[MUL.scala 105:13]
  assign m_111_io_x1 = r_282; // @[MUL.scala 103:13]
  assign m_111_io_x2 = r_283; // @[MUL.scala 104:13]
  assign m_111_io_x3 = r_284; // @[MUL.scala 105:13]
  assign m_112_io_in_0 = r_285; // @[MUL.scala 125:16]
  assign m_112_io_in_1 = r_286; // @[MUL.scala 126:16]
  assign m_113_io_x1 = r_287; // @[MUL.scala 103:13]
  assign m_113_io_x2 = r_288; // @[MUL.scala 104:13]
  assign m_113_io_x3 = r_289; // @[MUL.scala 105:13]
  assign m_114_io_x1 = r_290; // @[MUL.scala 103:13]
  assign m_114_io_x2 = r_291; // @[MUL.scala 104:13]
  assign m_114_io_x3 = r_292; // @[MUL.scala 105:13]
  assign m_115_io_x1 = r_293; // @[MUL.scala 103:13]
  assign m_115_io_x2 = r_294; // @[MUL.scala 104:13]
  assign m_115_io_x3 = r_295; // @[MUL.scala 105:13]
  assign m_116_io_x1 = r_296; // @[MUL.scala 103:13]
  assign m_116_io_x2 = r_297; // @[MUL.scala 104:13]
  assign m_116_io_x3 = r_298; // @[MUL.scala 105:13]
  assign m_117_io_x1 = r_299; // @[MUL.scala 103:13]
  assign m_117_io_x2 = r_300; // @[MUL.scala 104:13]
  assign m_117_io_x3 = r_301; // @[MUL.scala 105:13]
  assign m_118_io_in_0 = r_302; // @[MUL.scala 125:16]
  assign m_118_io_in_1 = r_303; // @[MUL.scala 126:16]
  assign m_119_io_x1 = r_304; // @[MUL.scala 103:13]
  assign m_119_io_x2 = r_305; // @[MUL.scala 104:13]
  assign m_119_io_x3 = r_306; // @[MUL.scala 105:13]
  assign m_120_io_x1 = r_307; // @[MUL.scala 103:13]
  assign m_120_io_x2 = r_308; // @[MUL.scala 104:13]
  assign m_120_io_x3 = r_309; // @[MUL.scala 105:13]
  assign m_121_io_x1 = r_310; // @[MUL.scala 103:13]
  assign m_121_io_x2 = r_311; // @[MUL.scala 104:13]
  assign m_121_io_x3 = r_312; // @[MUL.scala 105:13]
  assign m_122_io_x1 = r_313; // @[MUL.scala 103:13]
  assign m_122_io_x2 = r_314; // @[MUL.scala 104:13]
  assign m_122_io_x3 = r_315; // @[MUL.scala 105:13]
  assign m_123_io_x1 = r_316; // @[MUL.scala 103:13]
  assign m_123_io_x2 = r_317; // @[MUL.scala 104:13]
  assign m_123_io_x3 = r_318; // @[MUL.scala 105:13]
  assign m_124_io_in_0 = r_319; // @[MUL.scala 125:16]
  assign m_124_io_in_1 = r_320; // @[MUL.scala 126:16]
  assign m_125_io_x1 = r_321; // @[MUL.scala 103:13]
  assign m_125_io_x2 = r_322; // @[MUL.scala 104:13]
  assign m_125_io_x3 = r_323; // @[MUL.scala 105:13]
  assign m_126_io_x1 = r_324; // @[MUL.scala 103:13]
  assign m_126_io_x2 = r_325; // @[MUL.scala 104:13]
  assign m_126_io_x3 = r_326; // @[MUL.scala 105:13]
  assign m_127_io_x1 = r_327; // @[MUL.scala 103:13]
  assign m_127_io_x2 = r_328; // @[MUL.scala 104:13]
  assign m_127_io_x3 = r_329; // @[MUL.scala 105:13]
  assign m_128_io_x1 = r_330; // @[MUL.scala 103:13]
  assign m_128_io_x2 = r_331; // @[MUL.scala 104:13]
  assign m_128_io_x3 = r_332; // @[MUL.scala 105:13]
  assign m_129_io_x1 = r_333; // @[MUL.scala 103:13]
  assign m_129_io_x2 = r_334; // @[MUL.scala 104:13]
  assign m_129_io_x3 = r_335; // @[MUL.scala 105:13]
  assign m_130_io_in_0 = r_336; // @[MUL.scala 125:16]
  assign m_130_io_in_1 = r_337; // @[MUL.scala 126:16]
  assign m_131_io_x1 = r_338; // @[MUL.scala 103:13]
  assign m_131_io_x2 = r_339; // @[MUL.scala 104:13]
  assign m_131_io_x3 = r_340; // @[MUL.scala 105:13]
  assign m_132_io_x1 = r_341; // @[MUL.scala 103:13]
  assign m_132_io_x2 = r_342; // @[MUL.scala 104:13]
  assign m_132_io_x3 = r_343; // @[MUL.scala 105:13]
  assign m_133_io_x1 = r_344; // @[MUL.scala 103:13]
  assign m_133_io_x2 = r_345; // @[MUL.scala 104:13]
  assign m_133_io_x3 = r_346; // @[MUL.scala 105:13]
  assign m_134_io_x1 = r_347; // @[MUL.scala 103:13]
  assign m_134_io_x2 = r_348; // @[MUL.scala 104:13]
  assign m_134_io_x3 = r_349; // @[MUL.scala 105:13]
  assign m_135_io_x1 = r_350; // @[MUL.scala 103:13]
  assign m_135_io_x2 = r_351; // @[MUL.scala 104:13]
  assign m_135_io_x3 = r_352; // @[MUL.scala 105:13]
  assign m_136_io_in_0 = r_353; // @[MUL.scala 125:16]
  assign m_136_io_in_1 = r_354; // @[MUL.scala 126:16]
  assign m_137_io_x1 = r_355; // @[MUL.scala 103:13]
  assign m_137_io_x2 = r_356; // @[MUL.scala 104:13]
  assign m_137_io_x3 = r_357; // @[MUL.scala 105:13]
  assign m_138_io_x1 = r_358; // @[MUL.scala 103:13]
  assign m_138_io_x2 = r_359; // @[MUL.scala 104:13]
  assign m_138_io_x3 = r_360; // @[MUL.scala 105:13]
  assign m_139_io_x1 = r_361; // @[MUL.scala 103:13]
  assign m_139_io_x2 = r_362; // @[MUL.scala 104:13]
  assign m_139_io_x3 = r_363; // @[MUL.scala 105:13]
  assign m_140_io_x1 = r_364; // @[MUL.scala 103:13]
  assign m_140_io_x2 = r_365; // @[MUL.scala 104:13]
  assign m_140_io_x3 = r_366; // @[MUL.scala 105:13]
  assign m_141_io_x1 = r_367; // @[MUL.scala 103:13]
  assign m_141_io_x2 = r_368; // @[MUL.scala 104:13]
  assign m_141_io_x3 = r_369; // @[MUL.scala 105:13]
  assign m_142_io_in_0 = r_370; // @[MUL.scala 125:16]
  assign m_142_io_in_1 = r_371; // @[MUL.scala 126:16]
  assign m_143_io_x1 = r_372; // @[MUL.scala 103:13]
  assign m_143_io_x2 = r_373; // @[MUL.scala 104:13]
  assign m_143_io_x3 = r_374; // @[MUL.scala 105:13]
  assign m_144_io_x1 = r_375; // @[MUL.scala 103:13]
  assign m_144_io_x2 = r_376; // @[MUL.scala 104:13]
  assign m_144_io_x3 = r_377; // @[MUL.scala 105:13]
  assign m_145_io_x1 = r_378; // @[MUL.scala 103:13]
  assign m_145_io_x2 = r_379; // @[MUL.scala 104:13]
  assign m_145_io_x3 = r_380; // @[MUL.scala 105:13]
  assign m_146_io_x1 = r_381; // @[MUL.scala 103:13]
  assign m_146_io_x2 = r_382; // @[MUL.scala 104:13]
  assign m_146_io_x3 = r_383; // @[MUL.scala 105:13]
  assign m_147_io_x1 = r_384; // @[MUL.scala 103:13]
  assign m_147_io_x2 = r_385; // @[MUL.scala 104:13]
  assign m_147_io_x3 = r_386; // @[MUL.scala 105:13]
  assign m_148_io_in_0 = r_387; // @[MUL.scala 125:16]
  assign m_148_io_in_1 = r_388; // @[MUL.scala 126:16]
  assign m_149_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_149_io_x2 = r_390; // @[MUL.scala 104:13]
  assign m_149_io_x3 = r_391; // @[MUL.scala 105:13]
  assign m_150_io_x1 = r_392; // @[MUL.scala 103:13]
  assign m_150_io_x2 = r_393; // @[MUL.scala 104:13]
  assign m_150_io_x3 = r_394; // @[MUL.scala 105:13]
  assign m_151_io_x1 = r_395; // @[MUL.scala 103:13]
  assign m_151_io_x2 = r_396; // @[MUL.scala 104:13]
  assign m_151_io_x3 = r_397; // @[MUL.scala 105:13]
  assign m_152_io_x1 = r_398; // @[MUL.scala 103:13]
  assign m_152_io_x2 = r_399; // @[MUL.scala 104:13]
  assign m_152_io_x3 = r_400; // @[MUL.scala 105:13]
  assign m_153_io_x1 = r_401; // @[MUL.scala 103:13]
  assign m_153_io_x2 = r_402; // @[MUL.scala 104:13]
  assign m_153_io_x3 = r_403; // @[MUL.scala 105:13]
  assign m_154_io_x1 = r_405; // @[MUL.scala 103:13]
  assign m_154_io_x2 = r_406; // @[MUL.scala 104:13]
  assign m_154_io_x3 = r_407; // @[MUL.scala 105:13]
  assign m_155_io_x1 = r_408; // @[MUL.scala 103:13]
  assign m_155_io_x2 = r_409; // @[MUL.scala 104:13]
  assign m_155_io_x3 = r_410; // @[MUL.scala 105:13]
  assign m_156_io_x1 = r_411; // @[MUL.scala 103:13]
  assign m_156_io_x2 = r_412; // @[MUL.scala 104:13]
  assign m_156_io_x3 = r_413; // @[MUL.scala 105:13]
  assign m_157_io_x1 = r_414; // @[MUL.scala 103:13]
  assign m_157_io_x2 = r_415; // @[MUL.scala 104:13]
  assign m_157_io_x3 = r_416; // @[MUL.scala 105:13]
  assign m_158_io_x1 = r_417; // @[MUL.scala 103:13]
  assign m_158_io_x2 = r_418; // @[MUL.scala 104:13]
  assign m_158_io_x3 = r_419; // @[MUL.scala 105:13]
  assign m_159_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_159_io_x2 = r_421; // @[MUL.scala 104:13]
  assign m_159_io_x3 = r_422; // @[MUL.scala 105:13]
  assign m_160_io_x1 = r_423; // @[MUL.scala 103:13]
  assign m_160_io_x2 = r_424; // @[MUL.scala 104:13]
  assign m_160_io_x3 = r_425; // @[MUL.scala 105:13]
  assign m_161_io_x1 = r_426; // @[MUL.scala 103:13]
  assign m_161_io_x2 = r_427; // @[MUL.scala 104:13]
  assign m_161_io_x3 = r_428; // @[MUL.scala 105:13]
  assign m_162_io_x1 = r_429; // @[MUL.scala 103:13]
  assign m_162_io_x2 = r_430; // @[MUL.scala 104:13]
  assign m_162_io_x3 = r_431; // @[MUL.scala 105:13]
  assign m_163_io_x1 = r_432; // @[MUL.scala 103:13]
  assign m_163_io_x2 = r_433; // @[MUL.scala 104:13]
  assign m_163_io_x3 = r_434; // @[MUL.scala 105:13]
  assign m_164_io_x1 = r_435; // @[MUL.scala 103:13]
  assign m_164_io_x2 = r_436; // @[MUL.scala 104:13]
  assign m_164_io_x3 = r_437; // @[MUL.scala 105:13]
  assign m_165_io_x1 = r_438; // @[MUL.scala 103:13]
  assign m_165_io_x2 = r_439; // @[MUL.scala 104:13]
  assign m_165_io_x3 = r_440; // @[MUL.scala 105:13]
  assign m_166_io_x1 = r_441; // @[MUL.scala 103:13]
  assign m_166_io_x2 = r_442; // @[MUL.scala 104:13]
  assign m_166_io_x3 = r_443; // @[MUL.scala 105:13]
  assign m_167_io_x1 = r_444; // @[MUL.scala 103:13]
  assign m_167_io_x2 = r_445; // @[MUL.scala 104:13]
  assign m_167_io_x3 = r_446; // @[MUL.scala 105:13]
  assign m_168_io_in_0 = r_447; // @[MUL.scala 125:16]
  assign m_168_io_in_1 = r_448; // @[MUL.scala 126:16]
  assign m_169_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_169_io_x2 = r_450; // @[MUL.scala 104:13]
  assign m_169_io_x3 = r_451; // @[MUL.scala 105:13]
  assign m_170_io_x1 = r_452; // @[MUL.scala 103:13]
  assign m_170_io_x2 = r_453; // @[MUL.scala 104:13]
  assign m_170_io_x3 = r_454; // @[MUL.scala 105:13]
  assign m_171_io_x1 = r_455; // @[MUL.scala 103:13]
  assign m_171_io_x2 = r_456; // @[MUL.scala 104:13]
  assign m_171_io_x3 = r_457; // @[MUL.scala 105:13]
  assign m_172_io_x1 = r_458; // @[MUL.scala 103:13]
  assign m_172_io_x2 = r_459; // @[MUL.scala 104:13]
  assign m_172_io_x3 = r_460; // @[MUL.scala 105:13]
  assign m_173_io_in_0 = r_461; // @[MUL.scala 125:16]
  assign m_173_io_in_1 = r_462; // @[MUL.scala 126:16]
  assign m_174_io_x1 = r_463; // @[MUL.scala 103:13]
  assign m_174_io_x2 = r_464; // @[MUL.scala 104:13]
  assign m_174_io_x3 = r_465; // @[MUL.scala 105:13]
  assign m_175_io_x1 = r_466; // @[MUL.scala 103:13]
  assign m_175_io_x2 = r_467; // @[MUL.scala 104:13]
  assign m_175_io_x3 = r_468; // @[MUL.scala 105:13]
  assign m_176_io_x1 = r_469; // @[MUL.scala 103:13]
  assign m_176_io_x2 = r_470; // @[MUL.scala 104:13]
  assign m_176_io_x3 = r_471; // @[MUL.scala 105:13]
  assign m_177_io_x1 = r_472; // @[MUL.scala 103:13]
  assign m_177_io_x2 = r_473; // @[MUL.scala 104:13]
  assign m_177_io_x3 = r_474; // @[MUL.scala 105:13]
  assign m_178_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_178_io_x2 = r_477; // @[MUL.scala 104:13]
  assign m_178_io_x3 = r_478; // @[MUL.scala 105:13]
  assign m_179_io_x1 = r_479; // @[MUL.scala 103:13]
  assign m_179_io_x2 = r_480; // @[MUL.scala 104:13]
  assign m_179_io_x3 = r_481; // @[MUL.scala 105:13]
  assign m_180_io_x1 = r_482; // @[MUL.scala 103:13]
  assign m_180_io_x2 = r_483; // @[MUL.scala 104:13]
  assign m_180_io_x3 = r_484; // @[MUL.scala 105:13]
  assign m_181_io_x1 = r_485; // @[MUL.scala 103:13]
  assign m_181_io_x2 = r_486; // @[MUL.scala 104:13]
  assign m_181_io_x3 = r_487; // @[MUL.scala 105:13]
  assign m_182_io_x1 = r_489; // @[MUL.scala 103:13]
  assign m_182_io_x2 = r_490; // @[MUL.scala 104:13]
  assign m_182_io_x3 = r_491; // @[MUL.scala 105:13]
  assign m_183_io_x1 = r_492; // @[MUL.scala 103:13]
  assign m_183_io_x2 = r_493; // @[MUL.scala 104:13]
  assign m_183_io_x3 = r_494; // @[MUL.scala 105:13]
  assign m_184_io_x1 = r_495; // @[MUL.scala 103:13]
  assign m_184_io_x2 = r_496; // @[MUL.scala 104:13]
  assign m_184_io_x3 = r_497; // @[MUL.scala 105:13]
  assign m_185_io_x1 = r_498; // @[MUL.scala 103:13]
  assign m_185_io_x2 = r_499; // @[MUL.scala 104:13]
  assign m_185_io_x3 = r_500; // @[MUL.scala 105:13]
  assign m_186_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_186_io_x2 = r_502; // @[MUL.scala 104:13]
  assign m_186_io_x3 = r_503; // @[MUL.scala 105:13]
  assign m_187_io_x1 = r_504; // @[MUL.scala 103:13]
  assign m_187_io_x2 = r_505; // @[MUL.scala 104:13]
  assign m_187_io_x3 = r_506; // @[MUL.scala 105:13]
  assign m_188_io_x1 = r_507; // @[MUL.scala 103:13]
  assign m_188_io_x2 = r_508; // @[MUL.scala 104:13]
  assign m_188_io_x3 = r_509; // @[MUL.scala 105:13]
  assign m_189_io_x1 = r_510; // @[MUL.scala 103:13]
  assign m_189_io_x2 = r_511; // @[MUL.scala 104:13]
  assign m_189_io_x3 = r_512; // @[MUL.scala 105:13]
  assign m_190_io_x1 = r_513; // @[MUL.scala 103:13]
  assign m_190_io_x2 = r_514; // @[MUL.scala 104:13]
  assign m_190_io_x3 = r_515; // @[MUL.scala 105:13]
  assign m_191_io_x1 = r_516; // @[MUL.scala 103:13]
  assign m_191_io_x2 = r_517; // @[MUL.scala 104:13]
  assign m_191_io_x3 = r_518; // @[MUL.scala 105:13]
  assign m_192_io_x1 = r_519; // @[MUL.scala 103:13]
  assign m_192_io_x2 = r_520; // @[MUL.scala 104:13]
  assign m_192_io_x3 = r_521; // @[MUL.scala 105:13]
  assign m_193_io_in_0 = r_522; // @[MUL.scala 125:16]
  assign m_193_io_in_1 = r_523; // @[MUL.scala 126:16]
  assign m_194_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_194_io_x2 = r_525; // @[MUL.scala 104:13]
  assign m_194_io_x3 = r_526; // @[MUL.scala 105:13]
  assign m_195_io_x1 = r_527; // @[MUL.scala 103:13]
  assign m_195_io_x2 = r_528; // @[MUL.scala 104:13]
  assign m_195_io_x3 = r_529; // @[MUL.scala 105:13]
  assign m_196_io_x1 = r_530; // @[MUL.scala 103:13]
  assign m_196_io_x2 = r_531; // @[MUL.scala 104:13]
  assign m_196_io_x3 = r_532; // @[MUL.scala 105:13]
  assign m_197_io_in_0 = r_533; // @[MUL.scala 125:16]
  assign m_197_io_in_1 = r_534; // @[MUL.scala 126:16]
  assign m_198_io_x1 = r_535; // @[MUL.scala 103:13]
  assign m_198_io_x2 = r_536; // @[MUL.scala 104:13]
  assign m_198_io_x3 = r_537; // @[MUL.scala 105:13]
  assign m_199_io_x1 = r_538; // @[MUL.scala 103:13]
  assign m_199_io_x2 = r_539; // @[MUL.scala 104:13]
  assign m_199_io_x3 = r_540; // @[MUL.scala 105:13]
  assign m_200_io_x1 = r_541; // @[MUL.scala 103:13]
  assign m_200_io_x2 = r_542; // @[MUL.scala 104:13]
  assign m_200_io_x3 = r_543; // @[MUL.scala 105:13]
  assign m_201_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_201_io_x2 = r_546; // @[MUL.scala 104:13]
  assign m_201_io_x3 = r_547; // @[MUL.scala 105:13]
  assign m_202_io_x1 = r_548; // @[MUL.scala 103:13]
  assign m_202_io_x2 = r_549; // @[MUL.scala 104:13]
  assign m_202_io_x3 = r_550; // @[MUL.scala 105:13]
  assign m_203_io_x1 = r_551; // @[MUL.scala 103:13]
  assign m_203_io_x2 = r_552; // @[MUL.scala 104:13]
  assign m_203_io_x3 = r_553; // @[MUL.scala 105:13]
  assign m_204_io_x1 = r_555; // @[MUL.scala 103:13]
  assign m_204_io_x2 = r_556; // @[MUL.scala 104:13]
  assign m_204_io_x3 = r_557; // @[MUL.scala 105:13]
  assign m_205_io_x1 = r_558; // @[MUL.scala 103:13]
  assign m_205_io_x2 = r_559; // @[MUL.scala 104:13]
  assign m_205_io_x3 = r_560; // @[MUL.scala 105:13]
  assign m_206_io_x1 = r_561; // @[MUL.scala 103:13]
  assign m_206_io_x2 = r_562; // @[MUL.scala 104:13]
  assign m_206_io_x3 = r_563; // @[MUL.scala 105:13]
  assign m_207_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_207_io_x2 = r_565; // @[MUL.scala 104:13]
  assign m_207_io_x3 = r_566; // @[MUL.scala 105:13]
  assign m_208_io_x1 = r_567; // @[MUL.scala 103:13]
  assign m_208_io_x2 = r_568; // @[MUL.scala 104:13]
  assign m_208_io_x3 = r_569; // @[MUL.scala 105:13]
  assign m_209_io_x1 = r_570; // @[MUL.scala 103:13]
  assign m_209_io_x2 = r_571; // @[MUL.scala 104:13]
  assign m_209_io_x3 = r_572; // @[MUL.scala 105:13]
  assign m_210_io_x1 = r_573; // @[MUL.scala 103:13]
  assign m_210_io_x2 = r_574; // @[MUL.scala 104:13]
  assign m_210_io_x3 = r_575; // @[MUL.scala 105:13]
  assign m_211_io_x1 = r_576; // @[MUL.scala 103:13]
  assign m_211_io_x2 = r_577; // @[MUL.scala 104:13]
  assign m_211_io_x3 = r_578; // @[MUL.scala 105:13]
  assign m_212_io_in_0 = r_579; // @[MUL.scala 125:16]
  assign m_212_io_in_1 = r_580; // @[MUL.scala 126:16]
  assign m_213_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_213_io_x2 = r_582; // @[MUL.scala 104:13]
  assign m_213_io_x3 = r_583; // @[MUL.scala 105:13]
  assign m_214_io_x1 = r_584; // @[MUL.scala 103:13]
  assign m_214_io_x2 = r_585; // @[MUL.scala 104:13]
  assign m_214_io_x3 = r_586; // @[MUL.scala 105:13]
  assign m_215_io_in_0 = r_587; // @[MUL.scala 125:16]
  assign m_215_io_in_1 = r_588; // @[MUL.scala 126:16]
  assign m_216_io_x1 = r_589; // @[MUL.scala 103:13]
  assign m_216_io_x2 = r_590; // @[MUL.scala 104:13]
  assign m_216_io_x3 = r_591; // @[MUL.scala 105:13]
  assign m_217_io_x1 = r_592; // @[MUL.scala 103:13]
  assign m_217_io_x2 = r_593; // @[MUL.scala 104:13]
  assign m_217_io_x3 = r_594; // @[MUL.scala 105:13]
  assign m_218_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_218_io_x2 = r_597; // @[MUL.scala 104:13]
  assign m_218_io_x3 = r_598; // @[MUL.scala 105:13]
  assign m_219_io_x1 = r_599; // @[MUL.scala 103:13]
  assign m_219_io_x2 = r_600; // @[MUL.scala 104:13]
  assign m_219_io_x3 = r_601; // @[MUL.scala 105:13]
  assign m_220_io_x1 = r_603; // @[MUL.scala 103:13]
  assign m_220_io_x2 = r_604; // @[MUL.scala 104:13]
  assign m_220_io_x3 = r_605; // @[MUL.scala 105:13]
  assign m_221_io_x1 = r_606; // @[MUL.scala 103:13]
  assign m_221_io_x2 = r_607; // @[MUL.scala 104:13]
  assign m_221_io_x3 = r_608; // @[MUL.scala 105:13]
  assign m_222_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_222_io_x2 = r_610; // @[MUL.scala 104:13]
  assign m_222_io_x3 = r_611; // @[MUL.scala 105:13]
  assign m_223_io_x1 = r_612; // @[MUL.scala 103:13]
  assign m_223_io_x2 = r_613; // @[MUL.scala 104:13]
  assign m_223_io_x3 = r_614; // @[MUL.scala 105:13]
  assign m_224_io_x1 = r_615; // @[MUL.scala 103:13]
  assign m_224_io_x2 = r_616; // @[MUL.scala 104:13]
  assign m_224_io_x3 = r_617; // @[MUL.scala 105:13]
  assign m_225_io_in_0 = r_618; // @[MUL.scala 125:16]
  assign m_225_io_in_1 = r_619; // @[MUL.scala 126:16]
  assign m_226_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_226_io_x2 = r_621; // @[MUL.scala 104:13]
  assign m_226_io_x3 = r_622; // @[MUL.scala 105:13]
  assign m_227_io_in_0 = r_623; // @[MUL.scala 125:16]
  assign m_227_io_in_1 = r_624; // @[MUL.scala 126:16]
  assign m_228_io_x1 = r_625; // @[MUL.scala 103:13]
  assign m_228_io_x2 = r_626; // @[MUL.scala 104:13]
  assign m_228_io_x3 = r_627; // @[MUL.scala 105:13]
  assign m_229_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_229_io_x2 = r_630; // @[MUL.scala 104:13]
  assign m_229_io_x3 = r_631; // @[MUL.scala 105:13]
  assign m_230_io_x1 = r_633; // @[MUL.scala 103:13]
  assign m_230_io_x2 = r_634; // @[MUL.scala 104:13]
  assign m_230_io_x3 = r_635; // @[MUL.scala 105:13]
  assign m_231_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_231_io_x2 = r_637; // @[MUL.scala 104:13]
  assign m_231_io_x3 = r_638; // @[MUL.scala 105:13]
  assign m_232_io_in_0 = r_639; // @[MUL.scala 125:16]
  assign m_232_io_in_1 = r_640; // @[MUL.scala 126:16]
  assign m_233_io_in_0 = 1'h1; // @[MUL.scala 125:16]
  assign m_233_io_in_1 = r_642; // @[MUL.scala 126:16]
  assign m_234_io_in_0 = m_18_io_out_0; // @[MUL.scala 125:16]
  assign m_234_io_in_1 = m_17_io_out_1; // @[MUL.scala 126:16]
  assign m_235_io_in_0 = m_19_io_s; // @[MUL.scala 262:21]
  assign m_235_io_in_1 = m_18_io_out_1; // @[MUL.scala 126:16]
  assign m_236_io_in_0 = m_20_io_s; // @[MUL.scala 262:21]
  assign m_236_io_in_1 = m_19_io_cout; // @[MUL.scala 263:22]
  assign m_237_io_x1 = m_21_io_s; // @[MUL.scala 262:21]
  assign m_237_io_x2 = m_20_io_cout; // @[MUL.scala 263:22]
  assign m_237_io_x3 = r_13; // @[MUL.scala 105:13]
  assign m_238_io_x1 = m_22_io_s; // @[MUL.scala 262:21]
  assign m_238_io_x2 = m_21_io_cout; // @[MUL.scala 263:22]
  assign m_238_io_x3 = r_17; // @[MUL.scala 105:13]
  assign m_239_io_x1 = m_23_io_s; // @[MUL.scala 262:21]
  assign m_239_io_x2 = m_22_io_cout; // @[MUL.scala 263:22]
  assign m_239_io_x3 = m_24_io_out_0; // @[MUL.scala 105:13]
  assign m_240_io_x1 = m_25_io_s; // @[MUL.scala 262:21]
  assign m_240_io_x2 = m_23_io_cout; // @[MUL.scala 263:22]
  assign m_240_io_x3 = m_26_io_out_0; // @[MUL.scala 105:13]
  assign m_241_io_x1 = m_27_io_s; // @[MUL.scala 262:21]
  assign m_241_io_x2 = m_25_io_cout; // @[MUL.scala 263:22]
  assign m_241_io_x3 = m_28_io_s; // @[MUL.scala 262:21]
  assign m_242_io_x1 = m_29_io_s; // @[MUL.scala 262:21]
  assign m_242_io_x2 = m_27_io_cout; // @[MUL.scala 263:22]
  assign m_242_io_x3 = m_30_io_s; // @[MUL.scala 262:21]
  assign m_243_io_x1 = m_31_io_s; // @[MUL.scala 262:21]
  assign m_243_io_x2 = m_29_io_cout; // @[MUL.scala 263:22]
  assign m_243_io_x3 = m_32_io_s; // @[MUL.scala 262:21]
  assign m_244_io_in_0 = m_30_io_cout; // @[MUL.scala 263:22]
  assign m_244_io_in_1 = r_46; // @[MUL.scala 126:16]
  assign m_245_io_x1 = m_33_io_s; // @[MUL.scala 262:21]
  assign m_245_io_x2 = m_31_io_cout; // @[MUL.scala 263:22]
  assign m_245_io_x3 = m_34_io_s; // @[MUL.scala 262:21]
  assign m_246_io_in_0 = m_32_io_cout; // @[MUL.scala 263:22]
  assign m_246_io_in_1 = r_53; // @[MUL.scala 126:16]
  assign m_247_io_x1 = m_35_io_s; // @[MUL.scala 262:21]
  assign m_247_io_x2 = m_33_io_cout; // @[MUL.scala 263:22]
  assign m_247_io_x3 = m_36_io_s; // @[MUL.scala 262:21]
  assign m_248_io_in_0 = m_34_io_cout; // @[MUL.scala 263:22]
  assign m_248_io_in_1 = m_37_io_out_0; // @[MUL.scala 126:16]
  assign m_249_io_x1 = m_38_io_s; // @[MUL.scala 262:21]
  assign m_249_io_x2 = m_35_io_cout; // @[MUL.scala 263:22]
  assign m_249_io_x3 = m_39_io_s; // @[MUL.scala 262:21]
  assign m_250_io_x1 = m_36_io_cout; // @[MUL.scala 263:22]
  assign m_250_io_x2 = m_40_io_out_0; // @[MUL.scala 104:13]
  assign m_250_io_x3 = m_37_io_out_1; // @[MUL.scala 105:13]
  assign m_251_io_x1 = m_41_io_s; // @[MUL.scala 262:21]
  assign m_251_io_x2 = m_38_io_cout; // @[MUL.scala 263:22]
  assign m_251_io_x3 = m_42_io_s; // @[MUL.scala 262:21]
  assign m_252_io_x1 = m_39_io_cout; // @[MUL.scala 263:22]
  assign m_252_io_x2 = m_43_io_s; // @[MUL.scala 262:21]
  assign m_252_io_x3 = m_40_io_out_1; // @[MUL.scala 105:13]
  assign m_253_io_x1 = m_44_io_s; // @[MUL.scala 262:21]
  assign m_253_io_x2 = m_41_io_cout; // @[MUL.scala 263:22]
  assign m_253_io_x3 = m_45_io_s; // @[MUL.scala 262:21]
  assign m_254_io_x1 = m_42_io_cout; // @[MUL.scala 263:22]
  assign m_254_io_x2 = m_46_io_s; // @[MUL.scala 262:21]
  assign m_254_io_x3 = m_43_io_cout; // @[MUL.scala 263:22]
  assign m_255_io_x1 = m_47_io_s; // @[MUL.scala 262:21]
  assign m_255_io_x2 = m_44_io_cout; // @[MUL.scala 263:22]
  assign m_255_io_x3 = m_48_io_s; // @[MUL.scala 262:21]
  assign m_256_io_x1 = m_45_io_cout; // @[MUL.scala 263:22]
  assign m_256_io_x2 = m_49_io_s; // @[MUL.scala 262:21]
  assign m_256_io_x3 = m_46_io_cout; // @[MUL.scala 263:22]
  assign m_257_io_x1 = m_50_io_s; // @[MUL.scala 262:21]
  assign m_257_io_x2 = m_47_io_cout; // @[MUL.scala 263:22]
  assign m_257_io_x3 = m_51_io_s; // @[MUL.scala 262:21]
  assign m_258_io_x1 = m_48_io_cout; // @[MUL.scala 263:22]
  assign m_258_io_x2 = m_52_io_s; // @[MUL.scala 262:21]
  assign m_258_io_x3 = m_49_io_cout; // @[MUL.scala 263:22]
  assign m_259_io_x1 = m_53_io_s; // @[MUL.scala 262:21]
  assign m_259_io_x2 = m_50_io_cout; // @[MUL.scala 263:22]
  assign m_259_io_x3 = m_54_io_s; // @[MUL.scala 262:21]
  assign m_260_io_x1 = m_51_io_cout; // @[MUL.scala 263:22]
  assign m_260_io_x2 = m_55_io_s; // @[MUL.scala 262:21]
  assign m_260_io_x3 = m_52_io_cout; // @[MUL.scala 263:22]
  assign m_261_io_x1 = m_57_io_s; // @[MUL.scala 262:21]
  assign m_261_io_x2 = m_53_io_cout; // @[MUL.scala 263:22]
  assign m_261_io_x3 = m_58_io_s; // @[MUL.scala 262:21]
  assign m_262_io_x1 = m_54_io_cout; // @[MUL.scala 263:22]
  assign m_262_io_x2 = m_59_io_s; // @[MUL.scala 262:21]
  assign m_262_io_x3 = m_55_io_cout; // @[MUL.scala 263:22]
  assign m_263_io_in_0 = m_60_io_out_0; // @[MUL.scala 125:16]
  assign m_263_io_in_1 = m_56_io_out_1; // @[MUL.scala 126:16]
  assign m_264_io_x1 = m_61_io_s; // @[MUL.scala 262:21]
  assign m_264_io_x2 = m_57_io_cout; // @[MUL.scala 263:22]
  assign m_264_io_x3 = m_62_io_s; // @[MUL.scala 262:21]
  assign m_265_io_x1 = m_58_io_cout; // @[MUL.scala 263:22]
  assign m_265_io_x2 = m_63_io_s; // @[MUL.scala 262:21]
  assign m_265_io_x3 = m_59_io_cout; // @[MUL.scala 263:22]
  assign m_266_io_in_0 = m_64_io_s; // @[MUL.scala 262:21]
  assign m_266_io_in_1 = m_60_io_out_1; // @[MUL.scala 126:16]
  assign m_267_io_x1 = m_65_io_s; // @[MUL.scala 262:21]
  assign m_267_io_x2 = m_61_io_cout; // @[MUL.scala 263:22]
  assign m_267_io_x3 = m_66_io_s; // @[MUL.scala 262:21]
  assign m_268_io_x1 = m_62_io_cout; // @[MUL.scala 263:22]
  assign m_268_io_x2 = m_67_io_s; // @[MUL.scala 262:21]
  assign m_268_io_x3 = m_63_io_cout; // @[MUL.scala 263:22]
  assign m_269_io_in_0 = m_68_io_s; // @[MUL.scala 262:21]
  assign m_269_io_in_1 = m_64_io_cout; // @[MUL.scala 263:22]
  assign m_270_io_x1 = m_69_io_s; // @[MUL.scala 262:21]
  assign m_270_io_x2 = m_65_io_cout; // @[MUL.scala 263:22]
  assign m_270_io_x3 = m_70_io_s; // @[MUL.scala 262:21]
  assign m_271_io_x1 = m_66_io_cout; // @[MUL.scala 263:22]
  assign m_271_io_x2 = m_71_io_s; // @[MUL.scala 262:21]
  assign m_271_io_x3 = m_67_io_cout; // @[MUL.scala 263:22]
  assign m_272_io_x1 = m_72_io_s; // @[MUL.scala 262:21]
  assign m_272_io_x2 = m_68_io_cout; // @[MUL.scala 263:22]
  assign m_272_io_x3 = r_166; // @[MUL.scala 105:13]
  assign m_273_io_x1 = m_73_io_s; // @[MUL.scala 262:21]
  assign m_273_io_x2 = m_69_io_cout; // @[MUL.scala 263:22]
  assign m_273_io_x3 = m_74_io_s; // @[MUL.scala 262:21]
  assign m_274_io_x1 = m_70_io_cout; // @[MUL.scala 263:22]
  assign m_274_io_x2 = m_75_io_s; // @[MUL.scala 262:21]
  assign m_274_io_x3 = m_71_io_cout; // @[MUL.scala 263:22]
  assign m_275_io_x1 = m_76_io_s; // @[MUL.scala 262:21]
  assign m_275_io_x2 = m_72_io_cout; // @[MUL.scala 263:22]
  assign m_275_io_x3 = r_179; // @[MUL.scala 105:13]
  assign m_276_io_x1 = m_77_io_s; // @[MUL.scala 262:21]
  assign m_276_io_x2 = m_73_io_cout; // @[MUL.scala 263:22]
  assign m_276_io_x3 = m_78_io_s; // @[MUL.scala 262:21]
  assign m_277_io_x1 = m_74_io_cout; // @[MUL.scala 263:22]
  assign m_277_io_x2 = m_79_io_s; // @[MUL.scala 262:21]
  assign m_277_io_x3 = m_75_io_cout; // @[MUL.scala 263:22]
  assign m_278_io_x1 = m_80_io_s; // @[MUL.scala 262:21]
  assign m_278_io_x2 = m_76_io_cout; // @[MUL.scala 263:22]
  assign m_278_io_x3 = m_81_io_out_0; // @[MUL.scala 105:13]
  assign m_279_io_x1 = m_82_io_s; // @[MUL.scala 262:21]
  assign m_279_io_x2 = m_77_io_cout; // @[MUL.scala 263:22]
  assign m_279_io_x3 = m_83_io_s; // @[MUL.scala 262:21]
  assign m_280_io_x1 = m_78_io_cout; // @[MUL.scala 263:22]
  assign m_280_io_x2 = m_84_io_s; // @[MUL.scala 262:21]
  assign m_280_io_x3 = m_79_io_cout; // @[MUL.scala 263:22]
  assign m_281_io_x1 = m_85_io_s; // @[MUL.scala 262:21]
  assign m_281_io_x2 = m_80_io_cout; // @[MUL.scala 263:22]
  assign m_281_io_x3 = m_86_io_out_0; // @[MUL.scala 105:13]
  assign m_282_io_x1 = m_87_io_s; // @[MUL.scala 262:21]
  assign m_282_io_x2 = m_82_io_cout; // @[MUL.scala 263:22]
  assign m_282_io_x3 = m_88_io_s; // @[MUL.scala 262:21]
  assign m_283_io_x1 = m_83_io_cout; // @[MUL.scala 263:22]
  assign m_283_io_x2 = m_89_io_s; // @[MUL.scala 262:21]
  assign m_283_io_x3 = m_84_io_cout; // @[MUL.scala 263:22]
  assign m_284_io_x1 = m_90_io_s; // @[MUL.scala 262:21]
  assign m_284_io_x2 = m_85_io_cout; // @[MUL.scala 263:22]
  assign m_284_io_x3 = m_91_io_s; // @[MUL.scala 262:21]
  assign m_285_io_x1 = m_92_io_s; // @[MUL.scala 262:21]
  assign m_285_io_x2 = m_87_io_cout; // @[MUL.scala 263:22]
  assign m_285_io_x3 = m_93_io_s; // @[MUL.scala 262:21]
  assign m_286_io_x1 = m_88_io_cout; // @[MUL.scala 263:22]
  assign m_286_io_x2 = m_94_io_s; // @[MUL.scala 262:21]
  assign m_286_io_x3 = m_89_io_cout; // @[MUL.scala 263:22]
  assign m_287_io_x1 = m_95_io_s; // @[MUL.scala 262:21]
  assign m_287_io_x2 = m_90_io_cout; // @[MUL.scala 263:22]
  assign m_287_io_x3 = m_96_io_s; // @[MUL.scala 262:21]
  assign m_288_io_x1 = m_97_io_s; // @[MUL.scala 262:21]
  assign m_288_io_x2 = m_92_io_cout; // @[MUL.scala 263:22]
  assign m_288_io_x3 = m_98_io_s; // @[MUL.scala 262:21]
  assign m_289_io_x1 = m_93_io_cout; // @[MUL.scala 263:22]
  assign m_289_io_x2 = m_99_io_s; // @[MUL.scala 262:21]
  assign m_289_io_x3 = m_94_io_cout; // @[MUL.scala 263:22]
  assign m_290_io_x1 = m_100_io_s; // @[MUL.scala 262:21]
  assign m_290_io_x2 = m_95_io_cout; // @[MUL.scala 263:22]
  assign m_290_io_x3 = m_101_io_s; // @[MUL.scala 262:21]
  assign m_291_io_in_0 = m_96_io_cout; // @[MUL.scala 263:22]
  assign m_291_io_in_1 = r_253; // @[MUL.scala 126:16]
  assign m_292_io_x1 = m_102_io_s; // @[MUL.scala 262:21]
  assign m_292_io_x2 = m_97_io_cout; // @[MUL.scala 263:22]
  assign m_292_io_x3 = m_103_io_s; // @[MUL.scala 262:21]
  assign m_293_io_x1 = m_98_io_cout; // @[MUL.scala 263:22]
  assign m_293_io_x2 = m_104_io_s; // @[MUL.scala 262:21]
  assign m_293_io_x3 = m_99_io_cout; // @[MUL.scala 263:22]
  assign m_294_io_x1 = m_105_io_s; // @[MUL.scala 262:21]
  assign m_294_io_x2 = m_100_io_cout; // @[MUL.scala 263:22]
  assign m_294_io_x3 = m_106_io_s; // @[MUL.scala 262:21]
  assign m_295_io_in_0 = m_101_io_cout; // @[MUL.scala 263:22]
  assign m_295_io_in_1 = r_269; // @[MUL.scala 126:16]
  assign m_296_io_x1 = m_107_io_s; // @[MUL.scala 262:21]
  assign m_296_io_x2 = m_102_io_cout; // @[MUL.scala 263:22]
  assign m_296_io_x3 = m_108_io_s; // @[MUL.scala 262:21]
  assign m_297_io_x1 = m_103_io_cout; // @[MUL.scala 263:22]
  assign m_297_io_x2 = m_109_io_s; // @[MUL.scala 262:21]
  assign m_297_io_x3 = m_104_io_cout; // @[MUL.scala 263:22]
  assign m_298_io_x1 = m_110_io_s; // @[MUL.scala 262:21]
  assign m_298_io_x2 = m_105_io_cout; // @[MUL.scala 263:22]
  assign m_298_io_x3 = m_111_io_s; // @[MUL.scala 262:21]
  assign m_299_io_in_0 = m_106_io_cout; // @[MUL.scala 263:22]
  assign m_299_io_in_1 = m_112_io_out_0; // @[MUL.scala 126:16]
  assign m_300_io_x1 = m_113_io_s; // @[MUL.scala 262:21]
  assign m_300_io_x2 = m_107_io_cout; // @[MUL.scala 263:22]
  assign m_300_io_x3 = m_114_io_s; // @[MUL.scala 262:21]
  assign m_301_io_x1 = m_108_io_cout; // @[MUL.scala 263:22]
  assign m_301_io_x2 = m_115_io_s; // @[MUL.scala 262:21]
  assign m_301_io_x3 = m_109_io_cout; // @[MUL.scala 263:22]
  assign m_302_io_x1 = m_116_io_s; // @[MUL.scala 262:21]
  assign m_302_io_x2 = m_110_io_cout; // @[MUL.scala 263:22]
  assign m_302_io_x3 = m_117_io_s; // @[MUL.scala 262:21]
  assign m_303_io_x1 = m_111_io_cout; // @[MUL.scala 263:22]
  assign m_303_io_x2 = m_118_io_out_0; // @[MUL.scala 104:13]
  assign m_303_io_x3 = m_112_io_out_1; // @[MUL.scala 105:13]
  assign m_304_io_x1 = m_119_io_s; // @[MUL.scala 262:21]
  assign m_304_io_x2 = m_113_io_cout; // @[MUL.scala 263:22]
  assign m_304_io_x3 = m_120_io_s; // @[MUL.scala 262:21]
  assign m_305_io_x1 = m_114_io_cout; // @[MUL.scala 263:22]
  assign m_305_io_x2 = m_121_io_s; // @[MUL.scala 262:21]
  assign m_305_io_x3 = m_115_io_cout; // @[MUL.scala 263:22]
  assign m_306_io_x1 = m_122_io_s; // @[MUL.scala 262:21]
  assign m_306_io_x2 = m_116_io_cout; // @[MUL.scala 263:22]
  assign m_306_io_x3 = m_123_io_s; // @[MUL.scala 262:21]
  assign m_307_io_x1 = m_117_io_cout; // @[MUL.scala 263:22]
  assign m_307_io_x2 = m_124_io_out_0; // @[MUL.scala 104:13]
  assign m_307_io_x3 = m_118_io_out_1; // @[MUL.scala 105:13]
  assign m_308_io_x1 = m_125_io_s; // @[MUL.scala 262:21]
  assign m_308_io_x2 = m_119_io_cout; // @[MUL.scala 263:22]
  assign m_308_io_x3 = m_126_io_s; // @[MUL.scala 262:21]
  assign m_309_io_x1 = m_120_io_cout; // @[MUL.scala 263:22]
  assign m_309_io_x2 = m_127_io_s; // @[MUL.scala 262:21]
  assign m_309_io_x3 = m_121_io_cout; // @[MUL.scala 263:22]
  assign m_310_io_x1 = m_128_io_s; // @[MUL.scala 262:21]
  assign m_310_io_x2 = m_122_io_cout; // @[MUL.scala 263:22]
  assign m_310_io_x3 = m_129_io_s; // @[MUL.scala 262:21]
  assign m_311_io_x1 = m_123_io_cout; // @[MUL.scala 263:22]
  assign m_311_io_x2 = m_130_io_out_0; // @[MUL.scala 104:13]
  assign m_311_io_x3 = m_124_io_out_1; // @[MUL.scala 105:13]
  assign m_312_io_x1 = m_131_io_s; // @[MUL.scala 262:21]
  assign m_312_io_x2 = m_125_io_cout; // @[MUL.scala 263:22]
  assign m_312_io_x3 = m_132_io_s; // @[MUL.scala 262:21]
  assign m_313_io_x1 = m_126_io_cout; // @[MUL.scala 263:22]
  assign m_313_io_x2 = m_133_io_s; // @[MUL.scala 262:21]
  assign m_313_io_x3 = m_127_io_cout; // @[MUL.scala 263:22]
  assign m_314_io_x1 = m_134_io_s; // @[MUL.scala 262:21]
  assign m_314_io_x2 = m_128_io_cout; // @[MUL.scala 263:22]
  assign m_314_io_x3 = m_135_io_s; // @[MUL.scala 262:21]
  assign m_315_io_x1 = m_129_io_cout; // @[MUL.scala 263:22]
  assign m_315_io_x2 = m_136_io_out_0; // @[MUL.scala 104:13]
  assign m_315_io_x3 = m_130_io_out_1; // @[MUL.scala 105:13]
  assign m_316_io_x1 = m_137_io_s; // @[MUL.scala 262:21]
  assign m_316_io_x2 = m_131_io_cout; // @[MUL.scala 263:22]
  assign m_316_io_x3 = m_138_io_s; // @[MUL.scala 262:21]
  assign m_317_io_x1 = m_132_io_cout; // @[MUL.scala 263:22]
  assign m_317_io_x2 = m_139_io_s; // @[MUL.scala 262:21]
  assign m_317_io_x3 = m_133_io_cout; // @[MUL.scala 263:22]
  assign m_318_io_x1 = m_140_io_s; // @[MUL.scala 262:21]
  assign m_318_io_x2 = m_134_io_cout; // @[MUL.scala 263:22]
  assign m_318_io_x3 = m_141_io_s; // @[MUL.scala 262:21]
  assign m_319_io_x1 = m_135_io_cout; // @[MUL.scala 263:22]
  assign m_319_io_x2 = m_142_io_out_0; // @[MUL.scala 104:13]
  assign m_319_io_x3 = m_136_io_out_1; // @[MUL.scala 105:13]
  assign m_320_io_x1 = m_143_io_s; // @[MUL.scala 262:21]
  assign m_320_io_x2 = m_137_io_cout; // @[MUL.scala 263:22]
  assign m_320_io_x3 = m_144_io_s; // @[MUL.scala 262:21]
  assign m_321_io_x1 = m_138_io_cout; // @[MUL.scala 263:22]
  assign m_321_io_x2 = m_145_io_s; // @[MUL.scala 262:21]
  assign m_321_io_x3 = m_139_io_cout; // @[MUL.scala 263:22]
  assign m_322_io_x1 = m_146_io_s; // @[MUL.scala 262:21]
  assign m_322_io_x2 = m_140_io_cout; // @[MUL.scala 263:22]
  assign m_322_io_x3 = m_147_io_s; // @[MUL.scala 262:21]
  assign m_323_io_x1 = m_141_io_cout; // @[MUL.scala 263:22]
  assign m_323_io_x2 = m_148_io_out_0; // @[MUL.scala 104:13]
  assign m_323_io_x3 = m_142_io_out_1; // @[MUL.scala 105:13]
  assign m_324_io_x1 = m_149_io_s; // @[MUL.scala 262:21]
  assign m_324_io_x2 = m_143_io_cout; // @[MUL.scala 263:22]
  assign m_324_io_x3 = m_150_io_s; // @[MUL.scala 262:21]
  assign m_325_io_x1 = m_144_io_cout; // @[MUL.scala 263:22]
  assign m_325_io_x2 = m_151_io_s; // @[MUL.scala 262:21]
  assign m_325_io_x3 = m_145_io_cout; // @[MUL.scala 263:22]
  assign m_326_io_x1 = m_152_io_s; // @[MUL.scala 262:21]
  assign m_326_io_x2 = m_146_io_cout; // @[MUL.scala 263:22]
  assign m_326_io_x3 = m_153_io_s; // @[MUL.scala 262:21]
  assign m_327_io_x1 = m_147_io_cout; // @[MUL.scala 263:22]
  assign m_327_io_x2 = r_404; // @[MUL.scala 104:13]
  assign m_327_io_x3 = m_148_io_out_1; // @[MUL.scala 105:13]
  assign m_328_io_x1 = m_154_io_s; // @[MUL.scala 262:21]
  assign m_328_io_x2 = m_149_io_cout; // @[MUL.scala 263:22]
  assign m_328_io_x3 = m_155_io_s; // @[MUL.scala 262:21]
  assign m_329_io_x1 = m_150_io_cout; // @[MUL.scala 263:22]
  assign m_329_io_x2 = m_156_io_s; // @[MUL.scala 262:21]
  assign m_329_io_x3 = m_151_io_cout; // @[MUL.scala 263:22]
  assign m_330_io_x1 = m_157_io_s; // @[MUL.scala 262:21]
  assign m_330_io_x2 = m_152_io_cout; // @[MUL.scala 263:22]
  assign m_330_io_x3 = m_158_io_s; // @[MUL.scala 262:21]
  assign m_331_io_x1 = m_159_io_s; // @[MUL.scala 262:21]
  assign m_331_io_x2 = m_154_io_cout; // @[MUL.scala 263:22]
  assign m_331_io_x3 = m_160_io_s; // @[MUL.scala 262:21]
  assign m_332_io_x1 = m_155_io_cout; // @[MUL.scala 263:22]
  assign m_332_io_x2 = m_161_io_s; // @[MUL.scala 262:21]
  assign m_332_io_x3 = m_156_io_cout; // @[MUL.scala 263:22]
  assign m_333_io_x1 = m_162_io_s; // @[MUL.scala 262:21]
  assign m_333_io_x2 = m_157_io_cout; // @[MUL.scala 263:22]
  assign m_333_io_x3 = m_163_io_s; // @[MUL.scala 262:21]
  assign m_334_io_x1 = m_164_io_s; // @[MUL.scala 262:21]
  assign m_334_io_x2 = m_159_io_cout; // @[MUL.scala 263:22]
  assign m_334_io_x3 = m_165_io_s; // @[MUL.scala 262:21]
  assign m_335_io_x1 = m_160_io_cout; // @[MUL.scala 263:22]
  assign m_335_io_x2 = m_166_io_s; // @[MUL.scala 262:21]
  assign m_335_io_x3 = m_161_io_cout; // @[MUL.scala 263:22]
  assign m_336_io_x1 = m_167_io_s; // @[MUL.scala 262:21]
  assign m_336_io_x2 = m_162_io_cout; // @[MUL.scala 263:22]
  assign m_336_io_x3 = m_168_io_out_0; // @[MUL.scala 105:13]
  assign m_337_io_x1 = m_169_io_s; // @[MUL.scala 262:21]
  assign m_337_io_x2 = m_164_io_cout; // @[MUL.scala 263:22]
  assign m_337_io_x3 = m_170_io_s; // @[MUL.scala 262:21]
  assign m_338_io_x1 = m_165_io_cout; // @[MUL.scala 263:22]
  assign m_338_io_x2 = m_171_io_s; // @[MUL.scala 262:21]
  assign m_338_io_x3 = m_166_io_cout; // @[MUL.scala 263:22]
  assign m_339_io_x1 = m_172_io_s; // @[MUL.scala 262:21]
  assign m_339_io_x2 = m_167_io_cout; // @[MUL.scala 263:22]
  assign m_339_io_x3 = m_173_io_out_0; // @[MUL.scala 105:13]
  assign m_340_io_x1 = m_174_io_s; // @[MUL.scala 262:21]
  assign m_340_io_x2 = m_169_io_cout; // @[MUL.scala 263:22]
  assign m_340_io_x3 = m_175_io_s; // @[MUL.scala 262:21]
  assign m_341_io_x1 = m_170_io_cout; // @[MUL.scala 263:22]
  assign m_341_io_x2 = m_176_io_s; // @[MUL.scala 262:21]
  assign m_341_io_x3 = m_171_io_cout; // @[MUL.scala 263:22]
  assign m_342_io_x1 = m_177_io_s; // @[MUL.scala 262:21]
  assign m_342_io_x2 = m_172_io_cout; // @[MUL.scala 263:22]
  assign m_342_io_x3 = r_475; // @[MUL.scala 105:13]
  assign m_343_io_x1 = m_178_io_s; // @[MUL.scala 262:21]
  assign m_343_io_x2 = m_174_io_cout; // @[MUL.scala 263:22]
  assign m_343_io_x3 = m_179_io_s; // @[MUL.scala 262:21]
  assign m_344_io_x1 = m_175_io_cout; // @[MUL.scala 263:22]
  assign m_344_io_x2 = m_180_io_s; // @[MUL.scala 262:21]
  assign m_344_io_x3 = m_176_io_cout; // @[MUL.scala 263:22]
  assign m_345_io_x1 = m_181_io_s; // @[MUL.scala 262:21]
  assign m_345_io_x2 = m_177_io_cout; // @[MUL.scala 263:22]
  assign m_345_io_x3 = r_488; // @[MUL.scala 105:13]
  assign m_346_io_x1 = m_182_io_s; // @[MUL.scala 262:21]
  assign m_346_io_x2 = m_178_io_cout; // @[MUL.scala 263:22]
  assign m_346_io_x3 = m_183_io_s; // @[MUL.scala 262:21]
  assign m_347_io_x1 = m_179_io_cout; // @[MUL.scala 263:22]
  assign m_347_io_x2 = m_184_io_s; // @[MUL.scala 262:21]
  assign m_347_io_x3 = m_180_io_cout; // @[MUL.scala 263:22]
  assign m_348_io_in_0 = m_185_io_s; // @[MUL.scala 262:21]
  assign m_348_io_in_1 = m_181_io_cout; // @[MUL.scala 263:22]
  assign m_349_io_x1 = m_186_io_s; // @[MUL.scala 262:21]
  assign m_349_io_x2 = m_182_io_cout; // @[MUL.scala 263:22]
  assign m_349_io_x3 = m_187_io_s; // @[MUL.scala 262:21]
  assign m_350_io_x1 = m_183_io_cout; // @[MUL.scala 263:22]
  assign m_350_io_x2 = m_188_io_s; // @[MUL.scala 262:21]
  assign m_350_io_x3 = m_184_io_cout; // @[MUL.scala 263:22]
  assign m_351_io_in_0 = m_189_io_s; // @[MUL.scala 262:21]
  assign m_351_io_in_1 = m_185_io_cout; // @[MUL.scala 263:22]
  assign m_352_io_x1 = m_190_io_s; // @[MUL.scala 262:21]
  assign m_352_io_x2 = m_186_io_cout; // @[MUL.scala 263:22]
  assign m_352_io_x3 = m_191_io_s; // @[MUL.scala 262:21]
  assign m_353_io_x1 = m_187_io_cout; // @[MUL.scala 263:22]
  assign m_353_io_x2 = m_192_io_s; // @[MUL.scala 262:21]
  assign m_353_io_x3 = m_188_io_cout; // @[MUL.scala 263:22]
  assign m_354_io_in_0 = m_193_io_out_0; // @[MUL.scala 125:16]
  assign m_354_io_in_1 = m_189_io_cout; // @[MUL.scala 263:22]
  assign m_355_io_x1 = m_194_io_s; // @[MUL.scala 262:21]
  assign m_355_io_x2 = m_190_io_cout; // @[MUL.scala 263:22]
  assign m_355_io_x3 = m_195_io_s; // @[MUL.scala 262:21]
  assign m_356_io_x1 = m_191_io_cout; // @[MUL.scala 263:22]
  assign m_356_io_x2 = m_196_io_s; // @[MUL.scala 262:21]
  assign m_356_io_x3 = m_192_io_cout; // @[MUL.scala 263:22]
  assign m_357_io_in_0 = m_197_io_out_0; // @[MUL.scala 125:16]
  assign m_357_io_in_1 = m_193_io_out_1; // @[MUL.scala 126:16]
  assign m_358_io_x1 = m_198_io_s; // @[MUL.scala 262:21]
  assign m_358_io_x2 = m_194_io_cout; // @[MUL.scala 263:22]
  assign m_358_io_x3 = m_199_io_s; // @[MUL.scala 262:21]
  assign m_359_io_x1 = m_195_io_cout; // @[MUL.scala 263:22]
  assign m_359_io_x2 = m_200_io_s; // @[MUL.scala 262:21]
  assign m_359_io_x3 = m_196_io_cout; // @[MUL.scala 263:22]
  assign m_360_io_in_0 = r_544; // @[MUL.scala 125:16]
  assign m_360_io_in_1 = m_197_io_out_1; // @[MUL.scala 126:16]
  assign m_361_io_x1 = m_201_io_s; // @[MUL.scala 262:21]
  assign m_361_io_x2 = m_198_io_cout; // @[MUL.scala 263:22]
  assign m_361_io_x3 = m_202_io_s; // @[MUL.scala 262:21]
  assign m_362_io_x1 = m_199_io_cout; // @[MUL.scala 263:22]
  assign m_362_io_x2 = m_203_io_s; // @[MUL.scala 262:21]
  assign m_362_io_x3 = m_200_io_cout; // @[MUL.scala 263:22]
  assign m_363_io_x1 = m_204_io_s; // @[MUL.scala 262:21]
  assign m_363_io_x2 = m_201_io_cout; // @[MUL.scala 263:22]
  assign m_363_io_x3 = m_205_io_s; // @[MUL.scala 262:21]
  assign m_364_io_x1 = m_202_io_cout; // @[MUL.scala 263:22]
  assign m_364_io_x2 = m_206_io_s; // @[MUL.scala 262:21]
  assign m_364_io_x3 = m_203_io_cout; // @[MUL.scala 263:22]
  assign m_365_io_x1 = m_207_io_s; // @[MUL.scala 262:21]
  assign m_365_io_x2 = m_204_io_cout; // @[MUL.scala 263:22]
  assign m_365_io_x3 = m_208_io_s; // @[MUL.scala 262:21]
  assign m_366_io_x1 = m_205_io_cout; // @[MUL.scala 263:22]
  assign m_366_io_x2 = m_209_io_s; // @[MUL.scala 262:21]
  assign m_366_io_x3 = m_206_io_cout; // @[MUL.scala 263:22]
  assign m_367_io_x1 = m_210_io_s; // @[MUL.scala 262:21]
  assign m_367_io_x2 = m_207_io_cout; // @[MUL.scala 263:22]
  assign m_367_io_x3 = m_211_io_s; // @[MUL.scala 262:21]
  assign m_368_io_x1 = m_208_io_cout; // @[MUL.scala 263:22]
  assign m_368_io_x2 = m_212_io_out_0; // @[MUL.scala 104:13]
  assign m_368_io_x3 = m_209_io_cout; // @[MUL.scala 263:22]
  assign m_369_io_x1 = m_213_io_s; // @[MUL.scala 262:21]
  assign m_369_io_x2 = m_210_io_cout; // @[MUL.scala 263:22]
  assign m_369_io_x3 = m_214_io_s; // @[MUL.scala 262:21]
  assign m_370_io_x1 = m_211_io_cout; // @[MUL.scala 263:22]
  assign m_370_io_x2 = m_215_io_out_0; // @[MUL.scala 104:13]
  assign m_370_io_x3 = m_212_io_out_1; // @[MUL.scala 105:13]
  assign m_371_io_x1 = m_216_io_s; // @[MUL.scala 262:21]
  assign m_371_io_x2 = m_213_io_cout; // @[MUL.scala 263:22]
  assign m_371_io_x3 = m_217_io_s; // @[MUL.scala 262:21]
  assign m_372_io_x1 = m_214_io_cout; // @[MUL.scala 263:22]
  assign m_372_io_x2 = r_595; // @[MUL.scala 104:13]
  assign m_372_io_x3 = m_215_io_out_1; // @[MUL.scala 105:13]
  assign m_373_io_x1 = m_218_io_s; // @[MUL.scala 262:21]
  assign m_373_io_x2 = m_216_io_cout; // @[MUL.scala 263:22]
  assign m_373_io_x3 = m_219_io_s; // @[MUL.scala 262:21]
  assign m_374_io_in_0 = m_217_io_cout; // @[MUL.scala 263:22]
  assign m_374_io_in_1 = r_602; // @[MUL.scala 126:16]
  assign m_375_io_x1 = m_220_io_s; // @[MUL.scala 262:21]
  assign m_375_io_x2 = m_218_io_cout; // @[MUL.scala 263:22]
  assign m_375_io_x3 = m_221_io_s; // @[MUL.scala 262:21]
  assign m_376_io_x1 = m_222_io_s; // @[MUL.scala 262:21]
  assign m_376_io_x2 = m_220_io_cout; // @[MUL.scala 263:22]
  assign m_376_io_x3 = m_223_io_s; // @[MUL.scala 262:21]
  assign m_377_io_x1 = m_224_io_s; // @[MUL.scala 262:21]
  assign m_377_io_x2 = m_222_io_cout; // @[MUL.scala 263:22]
  assign m_377_io_x3 = m_225_io_out_0; // @[MUL.scala 105:13]
  assign m_378_io_x1 = m_226_io_s; // @[MUL.scala 262:21]
  assign m_378_io_x2 = m_224_io_cout; // @[MUL.scala 263:22]
  assign m_378_io_x3 = m_227_io_out_0; // @[MUL.scala 105:13]
  assign m_379_io_x1 = m_228_io_s; // @[MUL.scala 262:21]
  assign m_379_io_x2 = m_226_io_cout; // @[MUL.scala 263:22]
  assign m_379_io_x3 = r_628; // @[MUL.scala 105:13]
  assign m_380_io_x1 = m_229_io_s; // @[MUL.scala 262:21]
  assign m_380_io_x2 = m_228_io_cout; // @[MUL.scala 263:22]
  assign m_380_io_x3 = r_632; // @[MUL.scala 105:13]
  assign m_381_io_in_0 = m_230_io_s; // @[MUL.scala 262:21]
  assign m_381_io_in_1 = m_229_io_cout; // @[MUL.scala 263:22]
  assign m_382_io_in_0 = m_231_io_s; // @[MUL.scala 262:21]
  assign m_382_io_in_1 = m_230_io_cout; // @[MUL.scala 263:22]
  assign m_383_io_in_0 = m_232_io_out_0; // @[MUL.scala 125:16]
  assign m_383_io_in_1 = m_231_io_cout; // @[MUL.scala 263:22]
  assign m_384_io_in_0 = m_233_io_out_0; // @[MUL.scala 125:16]
  assign m_384_io_in_1 = m_232_io_out_1; // @[MUL.scala 126:16]
  assign m_385_io_in_0 = r_643; // @[MUL.scala 125:16]
  assign m_385_io_in_1 = m_233_io_out_1; // @[MUL.scala 126:16]
  assign m_386_io_in_0 = m_235_io_out_0; // @[MUL.scala 125:16]
  assign m_386_io_in_1 = m_234_io_out_1; // @[MUL.scala 126:16]
  assign m_387_io_in_0 = m_236_io_out_0; // @[MUL.scala 125:16]
  assign m_387_io_in_1 = m_235_io_out_1; // @[MUL.scala 126:16]
  assign m_388_io_in_0 = m_237_io_s; // @[MUL.scala 262:21]
  assign m_388_io_in_1 = m_236_io_out_1; // @[MUL.scala 126:16]
  assign m_389_io_in_0 = m_238_io_s; // @[MUL.scala 262:21]
  assign m_389_io_in_1 = m_237_io_cout; // @[MUL.scala 263:22]
  assign m_390_io_in_0 = m_239_io_s; // @[MUL.scala 262:21]
  assign m_390_io_in_1 = m_238_io_cout; // @[MUL.scala 263:22]
  assign m_391_io_x1 = m_240_io_s; // @[MUL.scala 262:21]
  assign m_391_io_x2 = m_239_io_cout; // @[MUL.scala 263:22]
  assign m_391_io_x3 = m_24_io_out_1; // @[MUL.scala 105:13]
  assign m_392_io_x1 = m_241_io_s; // @[MUL.scala 262:21]
  assign m_392_io_x2 = m_240_io_cout; // @[MUL.scala 263:22]
  assign m_392_io_x3 = m_26_io_out_1; // @[MUL.scala 105:13]
  assign m_393_io_x1 = m_242_io_s; // @[MUL.scala 262:21]
  assign m_393_io_x2 = m_241_io_cout; // @[MUL.scala 263:22]
  assign m_393_io_x3 = m_28_io_cout; // @[MUL.scala 263:22]
  assign m_394_io_x1 = m_243_io_s; // @[MUL.scala 262:21]
  assign m_394_io_x2 = m_242_io_cout; // @[MUL.scala 263:22]
  assign m_394_io_x3 = m_244_io_out_0; // @[MUL.scala 105:13]
  assign m_395_io_x1 = m_245_io_s; // @[MUL.scala 262:21]
  assign m_395_io_x2 = m_243_io_cout; // @[MUL.scala 263:22]
  assign m_395_io_x3 = m_246_io_out_0; // @[MUL.scala 105:13]
  assign m_396_io_x1 = m_247_io_s; // @[MUL.scala 262:21]
  assign m_396_io_x2 = m_245_io_cout; // @[MUL.scala 263:22]
  assign m_396_io_x3 = m_248_io_out_0; // @[MUL.scala 105:13]
  assign m_397_io_x1 = m_249_io_s; // @[MUL.scala 262:21]
  assign m_397_io_x2 = m_247_io_cout; // @[MUL.scala 263:22]
  assign m_397_io_x3 = m_250_io_s; // @[MUL.scala 262:21]
  assign m_398_io_x1 = m_251_io_s; // @[MUL.scala 262:21]
  assign m_398_io_x2 = m_249_io_cout; // @[MUL.scala 263:22]
  assign m_398_io_x3 = m_252_io_s; // @[MUL.scala 262:21]
  assign m_399_io_x1 = m_253_io_s; // @[MUL.scala 262:21]
  assign m_399_io_x2 = m_251_io_cout; // @[MUL.scala 263:22]
  assign m_399_io_x3 = m_254_io_s; // @[MUL.scala 262:21]
  assign m_400_io_x1 = m_255_io_s; // @[MUL.scala 262:21]
  assign m_400_io_x2 = m_253_io_cout; // @[MUL.scala 263:22]
  assign m_400_io_x3 = m_256_io_s; // @[MUL.scala 262:21]
  assign m_401_io_in_0 = m_254_io_cout; // @[MUL.scala 263:22]
  assign m_401_io_in_1 = r_97; // @[MUL.scala 126:16]
  assign m_402_io_x1 = m_257_io_s; // @[MUL.scala 262:21]
  assign m_402_io_x2 = m_255_io_cout; // @[MUL.scala 263:22]
  assign m_402_io_x3 = m_258_io_s; // @[MUL.scala 262:21]
  assign m_403_io_in_0 = m_256_io_cout; // @[MUL.scala 263:22]
  assign m_403_io_in_1 = r_107; // @[MUL.scala 126:16]
  assign m_404_io_x1 = m_259_io_s; // @[MUL.scala 262:21]
  assign m_404_io_x2 = m_257_io_cout; // @[MUL.scala 263:22]
  assign m_404_io_x3 = m_260_io_s; // @[MUL.scala 262:21]
  assign m_405_io_in_0 = m_258_io_cout; // @[MUL.scala 263:22]
  assign m_405_io_in_1 = m_56_io_out_0; // @[MUL.scala 126:16]
  assign m_406_io_x1 = m_261_io_s; // @[MUL.scala 262:21]
  assign m_406_io_x2 = m_259_io_cout; // @[MUL.scala 263:22]
  assign m_406_io_x3 = m_262_io_s; // @[MUL.scala 262:21]
  assign m_407_io_in_0 = m_260_io_cout; // @[MUL.scala 263:22]
  assign m_407_io_in_1 = m_263_io_out_0; // @[MUL.scala 126:16]
  assign m_408_io_x1 = m_264_io_s; // @[MUL.scala 262:21]
  assign m_408_io_x2 = m_261_io_cout; // @[MUL.scala 263:22]
  assign m_408_io_x3 = m_265_io_s; // @[MUL.scala 262:21]
  assign m_409_io_x1 = m_262_io_cout; // @[MUL.scala 263:22]
  assign m_409_io_x2 = m_266_io_out_0; // @[MUL.scala 104:13]
  assign m_409_io_x3 = m_263_io_out_1; // @[MUL.scala 105:13]
  assign m_410_io_x1 = m_267_io_s; // @[MUL.scala 262:21]
  assign m_410_io_x2 = m_264_io_cout; // @[MUL.scala 263:22]
  assign m_410_io_x3 = m_268_io_s; // @[MUL.scala 262:21]
  assign m_411_io_x1 = m_265_io_cout; // @[MUL.scala 263:22]
  assign m_411_io_x2 = m_269_io_out_0; // @[MUL.scala 104:13]
  assign m_411_io_x3 = m_266_io_out_1; // @[MUL.scala 105:13]
  assign m_412_io_x1 = m_270_io_s; // @[MUL.scala 262:21]
  assign m_412_io_x2 = m_267_io_cout; // @[MUL.scala 263:22]
  assign m_412_io_x3 = m_271_io_s; // @[MUL.scala 262:21]
  assign m_413_io_x1 = m_268_io_cout; // @[MUL.scala 263:22]
  assign m_413_io_x2 = m_272_io_s; // @[MUL.scala 262:21]
  assign m_413_io_x3 = m_269_io_out_1; // @[MUL.scala 105:13]
  assign m_414_io_x1 = m_273_io_s; // @[MUL.scala 262:21]
  assign m_414_io_x2 = m_270_io_cout; // @[MUL.scala 263:22]
  assign m_414_io_x3 = m_274_io_s; // @[MUL.scala 262:21]
  assign m_415_io_x1 = m_271_io_cout; // @[MUL.scala 263:22]
  assign m_415_io_x2 = m_275_io_s; // @[MUL.scala 262:21]
  assign m_415_io_x3 = m_272_io_cout; // @[MUL.scala 263:22]
  assign m_416_io_x1 = m_276_io_s; // @[MUL.scala 262:21]
  assign m_416_io_x2 = m_273_io_cout; // @[MUL.scala 263:22]
  assign m_416_io_x3 = m_277_io_s; // @[MUL.scala 262:21]
  assign m_417_io_x1 = m_274_io_cout; // @[MUL.scala 263:22]
  assign m_417_io_x2 = m_278_io_s; // @[MUL.scala 262:21]
  assign m_417_io_x3 = m_275_io_cout; // @[MUL.scala 263:22]
  assign m_418_io_x1 = m_279_io_s; // @[MUL.scala 262:21]
  assign m_418_io_x2 = m_276_io_cout; // @[MUL.scala 263:22]
  assign m_418_io_x3 = m_280_io_s; // @[MUL.scala 262:21]
  assign m_419_io_x1 = m_277_io_cout; // @[MUL.scala 263:22]
  assign m_419_io_x2 = m_281_io_s; // @[MUL.scala 262:21]
  assign m_419_io_x3 = m_278_io_cout; // @[MUL.scala 263:22]
  assign m_420_io_x1 = m_282_io_s; // @[MUL.scala 262:21]
  assign m_420_io_x2 = m_279_io_cout; // @[MUL.scala 263:22]
  assign m_420_io_x3 = m_283_io_s; // @[MUL.scala 262:21]
  assign m_421_io_x1 = m_280_io_cout; // @[MUL.scala 263:22]
  assign m_421_io_x2 = m_284_io_s; // @[MUL.scala 262:21]
  assign m_421_io_x3 = m_281_io_cout; // @[MUL.scala 263:22]
  assign m_422_io_x1 = m_285_io_s; // @[MUL.scala 262:21]
  assign m_422_io_x2 = m_282_io_cout; // @[MUL.scala 263:22]
  assign m_422_io_x3 = m_286_io_s; // @[MUL.scala 262:21]
  assign m_423_io_x1 = m_283_io_cout; // @[MUL.scala 263:22]
  assign m_423_io_x2 = m_287_io_s; // @[MUL.scala 262:21]
  assign m_423_io_x3 = m_284_io_cout; // @[MUL.scala 263:22]
  assign m_424_io_x1 = m_288_io_s; // @[MUL.scala 262:21]
  assign m_424_io_x2 = m_285_io_cout; // @[MUL.scala 263:22]
  assign m_424_io_x3 = m_289_io_s; // @[MUL.scala 262:21]
  assign m_425_io_x1 = m_286_io_cout; // @[MUL.scala 263:22]
  assign m_425_io_x2 = m_290_io_s; // @[MUL.scala 262:21]
  assign m_425_io_x3 = m_287_io_cout; // @[MUL.scala 263:22]
  assign m_426_io_x1 = m_292_io_s; // @[MUL.scala 262:21]
  assign m_426_io_x2 = m_288_io_cout; // @[MUL.scala 263:22]
  assign m_426_io_x3 = m_293_io_s; // @[MUL.scala 262:21]
  assign m_427_io_x1 = m_289_io_cout; // @[MUL.scala 263:22]
  assign m_427_io_x2 = m_294_io_s; // @[MUL.scala 262:21]
  assign m_427_io_x3 = m_290_io_cout; // @[MUL.scala 263:22]
  assign m_428_io_in_0 = m_295_io_out_0; // @[MUL.scala 125:16]
  assign m_428_io_in_1 = m_291_io_out_1; // @[MUL.scala 126:16]
  assign m_429_io_x1 = m_296_io_s; // @[MUL.scala 262:21]
  assign m_429_io_x2 = m_292_io_cout; // @[MUL.scala 263:22]
  assign m_429_io_x3 = m_297_io_s; // @[MUL.scala 262:21]
  assign m_430_io_x1 = m_293_io_cout; // @[MUL.scala 263:22]
  assign m_430_io_x2 = m_298_io_s; // @[MUL.scala 262:21]
  assign m_430_io_x3 = m_294_io_cout; // @[MUL.scala 263:22]
  assign m_431_io_in_0 = m_299_io_out_0; // @[MUL.scala 125:16]
  assign m_431_io_in_1 = m_295_io_out_1; // @[MUL.scala 126:16]
  assign m_432_io_x1 = m_300_io_s; // @[MUL.scala 262:21]
  assign m_432_io_x2 = m_296_io_cout; // @[MUL.scala 263:22]
  assign m_432_io_x3 = m_301_io_s; // @[MUL.scala 262:21]
  assign m_433_io_x1 = m_297_io_cout; // @[MUL.scala 263:22]
  assign m_433_io_x2 = m_302_io_s; // @[MUL.scala 262:21]
  assign m_433_io_x3 = m_298_io_cout; // @[MUL.scala 263:22]
  assign m_434_io_in_0 = m_303_io_s; // @[MUL.scala 262:21]
  assign m_434_io_in_1 = m_299_io_out_1; // @[MUL.scala 126:16]
  assign m_435_io_x1 = m_304_io_s; // @[MUL.scala 262:21]
  assign m_435_io_x2 = m_300_io_cout; // @[MUL.scala 263:22]
  assign m_435_io_x3 = m_305_io_s; // @[MUL.scala 262:21]
  assign m_436_io_x1 = m_301_io_cout; // @[MUL.scala 263:22]
  assign m_436_io_x2 = m_306_io_s; // @[MUL.scala 262:21]
  assign m_436_io_x3 = m_302_io_cout; // @[MUL.scala 263:22]
  assign m_437_io_in_0 = m_307_io_s; // @[MUL.scala 262:21]
  assign m_437_io_in_1 = m_303_io_cout; // @[MUL.scala 263:22]
  assign m_438_io_x1 = m_308_io_s; // @[MUL.scala 262:21]
  assign m_438_io_x2 = m_304_io_cout; // @[MUL.scala 263:22]
  assign m_438_io_x3 = m_309_io_s; // @[MUL.scala 262:21]
  assign m_439_io_x1 = m_305_io_cout; // @[MUL.scala 263:22]
  assign m_439_io_x2 = m_310_io_s; // @[MUL.scala 262:21]
  assign m_439_io_x3 = m_306_io_cout; // @[MUL.scala 263:22]
  assign m_440_io_in_0 = m_311_io_s; // @[MUL.scala 262:21]
  assign m_440_io_in_1 = m_307_io_cout; // @[MUL.scala 263:22]
  assign m_441_io_x1 = m_312_io_s; // @[MUL.scala 262:21]
  assign m_441_io_x2 = m_308_io_cout; // @[MUL.scala 263:22]
  assign m_441_io_x3 = m_313_io_s; // @[MUL.scala 262:21]
  assign m_442_io_x1 = m_309_io_cout; // @[MUL.scala 263:22]
  assign m_442_io_x2 = m_314_io_s; // @[MUL.scala 262:21]
  assign m_442_io_x3 = m_310_io_cout; // @[MUL.scala 263:22]
  assign m_443_io_in_0 = m_315_io_s; // @[MUL.scala 262:21]
  assign m_443_io_in_1 = m_311_io_cout; // @[MUL.scala 263:22]
  assign m_444_io_x1 = m_316_io_s; // @[MUL.scala 262:21]
  assign m_444_io_x2 = m_312_io_cout; // @[MUL.scala 263:22]
  assign m_444_io_x3 = m_317_io_s; // @[MUL.scala 262:21]
  assign m_445_io_x1 = m_313_io_cout; // @[MUL.scala 263:22]
  assign m_445_io_x2 = m_318_io_s; // @[MUL.scala 262:21]
  assign m_445_io_x3 = m_314_io_cout; // @[MUL.scala 263:22]
  assign m_446_io_in_0 = m_319_io_s; // @[MUL.scala 262:21]
  assign m_446_io_in_1 = m_315_io_cout; // @[MUL.scala 263:22]
  assign m_447_io_x1 = m_320_io_s; // @[MUL.scala 262:21]
  assign m_447_io_x2 = m_316_io_cout; // @[MUL.scala 263:22]
  assign m_447_io_x3 = m_321_io_s; // @[MUL.scala 262:21]
  assign m_448_io_x1 = m_317_io_cout; // @[MUL.scala 263:22]
  assign m_448_io_x2 = m_322_io_s; // @[MUL.scala 262:21]
  assign m_448_io_x3 = m_318_io_cout; // @[MUL.scala 263:22]
  assign m_449_io_in_0 = m_323_io_s; // @[MUL.scala 262:21]
  assign m_449_io_in_1 = m_319_io_cout; // @[MUL.scala 263:22]
  assign m_450_io_x1 = m_324_io_s; // @[MUL.scala 262:21]
  assign m_450_io_x2 = m_320_io_cout; // @[MUL.scala 263:22]
  assign m_450_io_x3 = m_325_io_s; // @[MUL.scala 262:21]
  assign m_451_io_x1 = m_321_io_cout; // @[MUL.scala 263:22]
  assign m_451_io_x2 = m_326_io_s; // @[MUL.scala 262:21]
  assign m_451_io_x3 = m_322_io_cout; // @[MUL.scala 263:22]
  assign m_452_io_in_0 = m_327_io_s; // @[MUL.scala 262:21]
  assign m_452_io_in_1 = m_323_io_cout; // @[MUL.scala 263:22]
  assign m_453_io_x1 = m_328_io_s; // @[MUL.scala 262:21]
  assign m_453_io_x2 = m_324_io_cout; // @[MUL.scala 263:22]
  assign m_453_io_x3 = m_329_io_s; // @[MUL.scala 262:21]
  assign m_454_io_x1 = m_325_io_cout; // @[MUL.scala 263:22]
  assign m_454_io_x2 = m_330_io_s; // @[MUL.scala 262:21]
  assign m_454_io_x3 = m_326_io_cout; // @[MUL.scala 263:22]
  assign m_455_io_in_0 = m_153_io_cout; // @[MUL.scala 263:22]
  assign m_455_io_in_1 = m_327_io_cout; // @[MUL.scala 263:22]
  assign m_456_io_x1 = m_331_io_s; // @[MUL.scala 262:21]
  assign m_456_io_x2 = m_328_io_cout; // @[MUL.scala 263:22]
  assign m_456_io_x3 = m_332_io_s; // @[MUL.scala 262:21]
  assign m_457_io_x1 = m_329_io_cout; // @[MUL.scala 263:22]
  assign m_457_io_x2 = m_333_io_s; // @[MUL.scala 262:21]
  assign m_457_io_x3 = m_330_io_cout; // @[MUL.scala 263:22]
  assign m_458_io_x1 = m_334_io_s; // @[MUL.scala 262:21]
  assign m_458_io_x2 = m_331_io_cout; // @[MUL.scala 263:22]
  assign m_458_io_x3 = m_335_io_s; // @[MUL.scala 262:21]
  assign m_459_io_x1 = m_332_io_cout; // @[MUL.scala 263:22]
  assign m_459_io_x2 = m_336_io_s; // @[MUL.scala 262:21]
  assign m_459_io_x3 = m_333_io_cout; // @[MUL.scala 263:22]
  assign m_460_io_x1 = m_337_io_s; // @[MUL.scala 262:21]
  assign m_460_io_x2 = m_334_io_cout; // @[MUL.scala 263:22]
  assign m_460_io_x3 = m_338_io_s; // @[MUL.scala 262:21]
  assign m_461_io_x1 = m_335_io_cout; // @[MUL.scala 263:22]
  assign m_461_io_x2 = m_339_io_s; // @[MUL.scala 262:21]
  assign m_461_io_x3 = m_336_io_cout; // @[MUL.scala 263:22]
  assign m_462_io_x1 = m_340_io_s; // @[MUL.scala 262:21]
  assign m_462_io_x2 = m_337_io_cout; // @[MUL.scala 263:22]
  assign m_462_io_x3 = m_341_io_s; // @[MUL.scala 262:21]
  assign m_463_io_x1 = m_338_io_cout; // @[MUL.scala 263:22]
  assign m_463_io_x2 = m_342_io_s; // @[MUL.scala 262:21]
  assign m_463_io_x3 = m_339_io_cout; // @[MUL.scala 263:22]
  assign m_464_io_x1 = m_343_io_s; // @[MUL.scala 262:21]
  assign m_464_io_x2 = m_340_io_cout; // @[MUL.scala 263:22]
  assign m_464_io_x3 = m_344_io_s; // @[MUL.scala 262:21]
  assign m_465_io_x1 = m_341_io_cout; // @[MUL.scala 263:22]
  assign m_465_io_x2 = m_345_io_s; // @[MUL.scala 262:21]
  assign m_465_io_x3 = m_342_io_cout; // @[MUL.scala 263:22]
  assign m_466_io_x1 = m_346_io_s; // @[MUL.scala 262:21]
  assign m_466_io_x2 = m_343_io_cout; // @[MUL.scala 263:22]
  assign m_466_io_x3 = m_347_io_s; // @[MUL.scala 262:21]
  assign m_467_io_x1 = m_344_io_cout; // @[MUL.scala 263:22]
  assign m_467_io_x2 = m_348_io_out_0; // @[MUL.scala 104:13]
  assign m_467_io_x3 = m_345_io_cout; // @[MUL.scala 263:22]
  assign m_468_io_x1 = m_349_io_s; // @[MUL.scala 262:21]
  assign m_468_io_x2 = m_346_io_cout; // @[MUL.scala 263:22]
  assign m_468_io_x3 = m_350_io_s; // @[MUL.scala 262:21]
  assign m_469_io_x1 = m_347_io_cout; // @[MUL.scala 263:22]
  assign m_469_io_x2 = m_351_io_out_0; // @[MUL.scala 104:13]
  assign m_469_io_x3 = m_348_io_out_1; // @[MUL.scala 105:13]
  assign m_470_io_x1 = m_352_io_s; // @[MUL.scala 262:21]
  assign m_470_io_x2 = m_349_io_cout; // @[MUL.scala 263:22]
  assign m_470_io_x3 = m_353_io_s; // @[MUL.scala 262:21]
  assign m_471_io_x1 = m_350_io_cout; // @[MUL.scala 263:22]
  assign m_471_io_x2 = m_354_io_out_0; // @[MUL.scala 104:13]
  assign m_471_io_x3 = m_351_io_out_1; // @[MUL.scala 105:13]
  assign m_472_io_x1 = m_355_io_s; // @[MUL.scala 262:21]
  assign m_472_io_x2 = m_352_io_cout; // @[MUL.scala 263:22]
  assign m_472_io_x3 = m_356_io_s; // @[MUL.scala 262:21]
  assign m_473_io_x1 = m_353_io_cout; // @[MUL.scala 263:22]
  assign m_473_io_x2 = m_357_io_out_0; // @[MUL.scala 104:13]
  assign m_473_io_x3 = m_354_io_out_1; // @[MUL.scala 105:13]
  assign m_474_io_x1 = m_358_io_s; // @[MUL.scala 262:21]
  assign m_474_io_x2 = m_355_io_cout; // @[MUL.scala 263:22]
  assign m_474_io_x3 = m_359_io_s; // @[MUL.scala 262:21]
  assign m_475_io_x1 = m_356_io_cout; // @[MUL.scala 263:22]
  assign m_475_io_x2 = m_360_io_out_0; // @[MUL.scala 104:13]
  assign m_475_io_x3 = m_357_io_out_1; // @[MUL.scala 105:13]
  assign m_476_io_x1 = m_361_io_s; // @[MUL.scala 262:21]
  assign m_476_io_x2 = m_358_io_cout; // @[MUL.scala 263:22]
  assign m_476_io_x3 = m_362_io_s; // @[MUL.scala 262:21]
  assign m_477_io_x1 = m_359_io_cout; // @[MUL.scala 263:22]
  assign m_477_io_x2 = r_554; // @[MUL.scala 104:13]
  assign m_477_io_x3 = m_360_io_out_1; // @[MUL.scala 105:13]
  assign m_478_io_x1 = m_363_io_s; // @[MUL.scala 262:21]
  assign m_478_io_x2 = m_361_io_cout; // @[MUL.scala 263:22]
  assign m_478_io_x3 = m_364_io_s; // @[MUL.scala 262:21]
  assign m_479_io_x1 = m_365_io_s; // @[MUL.scala 262:21]
  assign m_479_io_x2 = m_363_io_cout; // @[MUL.scala 263:22]
  assign m_479_io_x3 = m_366_io_s; // @[MUL.scala 262:21]
  assign m_480_io_x1 = m_367_io_s; // @[MUL.scala 262:21]
  assign m_480_io_x2 = m_365_io_cout; // @[MUL.scala 263:22]
  assign m_480_io_x3 = m_368_io_s; // @[MUL.scala 262:21]
  assign m_481_io_x1 = m_369_io_s; // @[MUL.scala 262:21]
  assign m_481_io_x2 = m_367_io_cout; // @[MUL.scala 263:22]
  assign m_481_io_x3 = m_370_io_s; // @[MUL.scala 262:21]
  assign m_482_io_x1 = m_371_io_s; // @[MUL.scala 262:21]
  assign m_482_io_x2 = m_369_io_cout; // @[MUL.scala 263:22]
  assign m_482_io_x3 = m_372_io_s; // @[MUL.scala 262:21]
  assign m_483_io_x1 = m_373_io_s; // @[MUL.scala 262:21]
  assign m_483_io_x2 = m_371_io_cout; // @[MUL.scala 263:22]
  assign m_483_io_x3 = m_374_io_out_0; // @[MUL.scala 105:13]
  assign m_484_io_x1 = m_375_io_s; // @[MUL.scala 262:21]
  assign m_484_io_x2 = m_373_io_cout; // @[MUL.scala 263:22]
  assign m_484_io_x3 = m_219_io_cout; // @[MUL.scala 263:22]
  assign m_485_io_x1 = m_376_io_s; // @[MUL.scala 262:21]
  assign m_485_io_x2 = m_375_io_cout; // @[MUL.scala 263:22]
  assign m_485_io_x3 = m_221_io_cout; // @[MUL.scala 263:22]
  assign m_486_io_x1 = m_377_io_s; // @[MUL.scala 262:21]
  assign m_486_io_x2 = m_376_io_cout; // @[MUL.scala 263:22]
  assign m_486_io_x3 = m_223_io_cout; // @[MUL.scala 263:22]
  assign m_487_io_x1 = m_378_io_s; // @[MUL.scala 262:21]
  assign m_487_io_x2 = m_377_io_cout; // @[MUL.scala 263:22]
  assign m_487_io_x3 = m_225_io_out_1; // @[MUL.scala 105:13]
  assign m_488_io_x1 = m_379_io_s; // @[MUL.scala 262:21]
  assign m_488_io_x2 = m_378_io_cout; // @[MUL.scala 263:22]
  assign m_488_io_x3 = m_227_io_out_1; // @[MUL.scala 105:13]
  assign m_489_io_in_0 = m_380_io_s; // @[MUL.scala 262:21]
  assign m_489_io_in_1 = m_379_io_cout; // @[MUL.scala 263:22]
  assign m_490_io_in_0 = m_381_io_out_0; // @[MUL.scala 125:16]
  assign m_490_io_in_1 = m_380_io_cout; // @[MUL.scala 263:22]
  assign m_491_io_in_0 = m_382_io_out_0; // @[MUL.scala 125:16]
  assign m_491_io_in_1 = m_381_io_out_1; // @[MUL.scala 126:16]
  assign m_492_io_in_0 = m_383_io_out_0; // @[MUL.scala 125:16]
  assign m_492_io_in_1 = m_382_io_out_1; // @[MUL.scala 126:16]
  assign m_493_io_in_0 = m_384_io_out_0; // @[MUL.scala 125:16]
  assign m_493_io_in_1 = m_383_io_out_1; // @[MUL.scala 126:16]
  assign m_494_io_in_0 = m_385_io_out_0; // @[MUL.scala 125:16]
  assign m_494_io_in_1 = m_384_io_out_1; // @[MUL.scala 126:16]
  assign m_495_io_in_0 = m_387_io_out_0; // @[MUL.scala 125:16]
  assign m_495_io_in_1 = m_386_io_out_1; // @[MUL.scala 126:16]
  assign m_496_io_in_0 = m_388_io_out_0; // @[MUL.scala 125:16]
  assign m_496_io_in_1 = m_387_io_out_1; // @[MUL.scala 126:16]
  assign m_497_io_in_0 = m_389_io_out_0; // @[MUL.scala 125:16]
  assign m_497_io_in_1 = m_388_io_out_1; // @[MUL.scala 126:16]
  assign m_498_io_in_0 = m_390_io_out_0; // @[MUL.scala 125:16]
  assign m_498_io_in_1 = m_389_io_out_1; // @[MUL.scala 126:16]
  assign m_499_io_in_0 = m_391_io_s; // @[MUL.scala 262:21]
  assign m_499_io_in_1 = m_390_io_out_1; // @[MUL.scala 126:16]
  assign m_500_io_in_0 = m_392_io_s; // @[MUL.scala 262:21]
  assign m_500_io_in_1 = m_391_io_cout; // @[MUL.scala 263:22]
  assign m_501_io_in_0 = m_393_io_s; // @[MUL.scala 262:21]
  assign m_501_io_in_1 = m_392_io_cout; // @[MUL.scala 263:22]
  assign m_502_io_in_0 = m_394_io_s; // @[MUL.scala 262:21]
  assign m_502_io_in_1 = m_393_io_cout; // @[MUL.scala 263:22]
  assign m_503_io_x1 = m_395_io_s; // @[MUL.scala 262:21]
  assign m_503_io_x2 = m_394_io_cout; // @[MUL.scala 263:22]
  assign m_503_io_x3 = m_244_io_out_1; // @[MUL.scala 105:13]
  assign m_504_io_x1 = m_396_io_s; // @[MUL.scala 262:21]
  assign m_504_io_x2 = m_395_io_cout; // @[MUL.scala 263:22]
  assign m_504_io_x3 = m_246_io_out_1; // @[MUL.scala 105:13]
  assign m_505_io_x1 = m_397_io_s; // @[MUL.scala 262:21]
  assign m_505_io_x2 = m_396_io_cout; // @[MUL.scala 263:22]
  assign m_505_io_x3 = m_248_io_out_1; // @[MUL.scala 105:13]
  assign m_506_io_x1 = m_398_io_s; // @[MUL.scala 262:21]
  assign m_506_io_x2 = m_397_io_cout; // @[MUL.scala 263:22]
  assign m_506_io_x3 = m_250_io_cout; // @[MUL.scala 263:22]
  assign m_507_io_x1 = m_399_io_s; // @[MUL.scala 262:21]
  assign m_507_io_x2 = m_398_io_cout; // @[MUL.scala 263:22]
  assign m_507_io_x3 = m_252_io_cout; // @[MUL.scala 263:22]
  assign m_508_io_x1 = m_400_io_s; // @[MUL.scala 262:21]
  assign m_508_io_x2 = m_399_io_cout; // @[MUL.scala 263:22]
  assign m_508_io_x3 = m_401_io_out_0; // @[MUL.scala 105:13]
  assign m_509_io_x1 = m_402_io_s; // @[MUL.scala 262:21]
  assign m_509_io_x2 = m_400_io_cout; // @[MUL.scala 263:22]
  assign m_509_io_x3 = m_403_io_out_0; // @[MUL.scala 105:13]
  assign m_510_io_x1 = m_404_io_s; // @[MUL.scala 262:21]
  assign m_510_io_x2 = m_402_io_cout; // @[MUL.scala 263:22]
  assign m_510_io_x3 = m_405_io_out_0; // @[MUL.scala 105:13]
  assign m_511_io_x1 = m_406_io_s; // @[MUL.scala 262:21]
  assign m_511_io_x2 = m_404_io_cout; // @[MUL.scala 263:22]
  assign m_511_io_x3 = m_407_io_out_0; // @[MUL.scala 105:13]
  assign m_512_io_x1 = m_408_io_s; // @[MUL.scala 262:21]
  assign m_512_io_x2 = m_406_io_cout; // @[MUL.scala 263:22]
  assign m_512_io_x3 = m_409_io_s; // @[MUL.scala 262:21]
  assign m_513_io_x1 = m_410_io_s; // @[MUL.scala 262:21]
  assign m_513_io_x2 = m_408_io_cout; // @[MUL.scala 263:22]
  assign m_513_io_x3 = m_411_io_s; // @[MUL.scala 262:21]
  assign m_514_io_x1 = m_412_io_s; // @[MUL.scala 262:21]
  assign m_514_io_x2 = m_410_io_cout; // @[MUL.scala 263:22]
  assign m_514_io_x3 = m_413_io_s; // @[MUL.scala 262:21]
  assign m_515_io_x1 = m_414_io_s; // @[MUL.scala 262:21]
  assign m_515_io_x2 = m_412_io_cout; // @[MUL.scala 263:22]
  assign m_515_io_x3 = m_415_io_s; // @[MUL.scala 262:21]
  assign m_516_io_x1 = m_416_io_s; // @[MUL.scala 262:21]
  assign m_516_io_x2 = m_414_io_cout; // @[MUL.scala 263:22]
  assign m_516_io_x3 = m_417_io_s; // @[MUL.scala 262:21]
  assign m_517_io_x1 = m_418_io_s; // @[MUL.scala 262:21]
  assign m_517_io_x2 = m_416_io_cout; // @[MUL.scala 263:22]
  assign m_517_io_x3 = m_419_io_s; // @[MUL.scala 262:21]
  assign m_518_io_in_0 = m_417_io_cout; // @[MUL.scala 263:22]
  assign m_518_io_in_1 = m_81_io_out_1; // @[MUL.scala 126:16]
  assign m_519_io_x1 = m_420_io_s; // @[MUL.scala 262:21]
  assign m_519_io_x2 = m_418_io_cout; // @[MUL.scala 263:22]
  assign m_519_io_x3 = m_421_io_s; // @[MUL.scala 262:21]
  assign m_520_io_in_0 = m_419_io_cout; // @[MUL.scala 263:22]
  assign m_520_io_in_1 = m_86_io_out_1; // @[MUL.scala 126:16]
  assign m_521_io_x1 = m_422_io_s; // @[MUL.scala 262:21]
  assign m_521_io_x2 = m_420_io_cout; // @[MUL.scala 263:22]
  assign m_521_io_x3 = m_423_io_s; // @[MUL.scala 262:21]
  assign m_522_io_in_0 = m_421_io_cout; // @[MUL.scala 263:22]
  assign m_522_io_in_1 = m_91_io_cout; // @[MUL.scala 263:22]
  assign m_523_io_x1 = m_424_io_s; // @[MUL.scala 262:21]
  assign m_523_io_x2 = m_422_io_cout; // @[MUL.scala 263:22]
  assign m_523_io_x3 = m_425_io_s; // @[MUL.scala 262:21]
  assign m_524_io_in_0 = m_423_io_cout; // @[MUL.scala 263:22]
  assign m_524_io_in_1 = m_291_io_out_0; // @[MUL.scala 126:16]
  assign m_525_io_x1 = m_426_io_s; // @[MUL.scala 262:21]
  assign m_525_io_x2 = m_424_io_cout; // @[MUL.scala 263:22]
  assign m_525_io_x3 = m_427_io_s; // @[MUL.scala 262:21]
  assign m_526_io_in_0 = m_425_io_cout; // @[MUL.scala 263:22]
  assign m_526_io_in_1 = m_428_io_out_0; // @[MUL.scala 126:16]
  assign m_527_io_x1 = m_429_io_s; // @[MUL.scala 262:21]
  assign m_527_io_x2 = m_426_io_cout; // @[MUL.scala 263:22]
  assign m_527_io_x3 = m_430_io_s; // @[MUL.scala 262:21]
  assign m_528_io_x1 = m_427_io_cout; // @[MUL.scala 263:22]
  assign m_528_io_x2 = m_431_io_out_0; // @[MUL.scala 104:13]
  assign m_528_io_x3 = m_428_io_out_1; // @[MUL.scala 105:13]
  assign m_529_io_x1 = m_432_io_s; // @[MUL.scala 262:21]
  assign m_529_io_x2 = m_429_io_cout; // @[MUL.scala 263:22]
  assign m_529_io_x3 = m_433_io_s; // @[MUL.scala 262:21]
  assign m_530_io_x1 = m_430_io_cout; // @[MUL.scala 263:22]
  assign m_530_io_x2 = m_434_io_out_0; // @[MUL.scala 104:13]
  assign m_530_io_x3 = m_431_io_out_1; // @[MUL.scala 105:13]
  assign m_531_io_x1 = m_435_io_s; // @[MUL.scala 262:21]
  assign m_531_io_x2 = m_432_io_cout; // @[MUL.scala 263:22]
  assign m_531_io_x3 = m_436_io_s; // @[MUL.scala 262:21]
  assign m_532_io_x1 = m_433_io_cout; // @[MUL.scala 263:22]
  assign m_532_io_x2 = m_437_io_out_0; // @[MUL.scala 104:13]
  assign m_532_io_x3 = m_434_io_out_1; // @[MUL.scala 105:13]
  assign m_533_io_x1 = m_438_io_s; // @[MUL.scala 262:21]
  assign m_533_io_x2 = m_435_io_cout; // @[MUL.scala 263:22]
  assign m_533_io_x3 = m_439_io_s; // @[MUL.scala 262:21]
  assign m_534_io_x1 = m_436_io_cout; // @[MUL.scala 263:22]
  assign m_534_io_x2 = m_440_io_out_0; // @[MUL.scala 104:13]
  assign m_534_io_x3 = m_437_io_out_1; // @[MUL.scala 105:13]
  assign m_535_io_x1 = m_441_io_s; // @[MUL.scala 262:21]
  assign m_535_io_x2 = m_438_io_cout; // @[MUL.scala 263:22]
  assign m_535_io_x3 = m_442_io_s; // @[MUL.scala 262:21]
  assign m_536_io_x1 = m_439_io_cout; // @[MUL.scala 263:22]
  assign m_536_io_x2 = m_443_io_out_0; // @[MUL.scala 104:13]
  assign m_536_io_x3 = m_440_io_out_1; // @[MUL.scala 105:13]
  assign m_537_io_x1 = m_444_io_s; // @[MUL.scala 262:21]
  assign m_537_io_x2 = m_441_io_cout; // @[MUL.scala 263:22]
  assign m_537_io_x3 = m_445_io_s; // @[MUL.scala 262:21]
  assign m_538_io_x1 = m_442_io_cout; // @[MUL.scala 263:22]
  assign m_538_io_x2 = m_446_io_out_0; // @[MUL.scala 104:13]
  assign m_538_io_x3 = m_443_io_out_1; // @[MUL.scala 105:13]
  assign m_539_io_x1 = m_447_io_s; // @[MUL.scala 262:21]
  assign m_539_io_x2 = m_444_io_cout; // @[MUL.scala 263:22]
  assign m_539_io_x3 = m_448_io_s; // @[MUL.scala 262:21]
  assign m_540_io_x1 = m_445_io_cout; // @[MUL.scala 263:22]
  assign m_540_io_x2 = m_449_io_out_0; // @[MUL.scala 104:13]
  assign m_540_io_x3 = m_446_io_out_1; // @[MUL.scala 105:13]
  assign m_541_io_x1 = m_450_io_s; // @[MUL.scala 262:21]
  assign m_541_io_x2 = m_447_io_cout; // @[MUL.scala 263:22]
  assign m_541_io_x3 = m_451_io_s; // @[MUL.scala 262:21]
  assign m_542_io_x1 = m_448_io_cout; // @[MUL.scala 263:22]
  assign m_542_io_x2 = m_452_io_out_0; // @[MUL.scala 104:13]
  assign m_542_io_x3 = m_449_io_out_1; // @[MUL.scala 105:13]
  assign m_543_io_x1 = m_453_io_s; // @[MUL.scala 262:21]
  assign m_543_io_x2 = m_450_io_cout; // @[MUL.scala 263:22]
  assign m_543_io_x3 = m_454_io_s; // @[MUL.scala 262:21]
  assign m_544_io_x1 = m_451_io_cout; // @[MUL.scala 263:22]
  assign m_544_io_x2 = m_455_io_out_0; // @[MUL.scala 104:13]
  assign m_544_io_x3 = m_452_io_out_1; // @[MUL.scala 105:13]
  assign m_545_io_x1 = m_456_io_s; // @[MUL.scala 262:21]
  assign m_545_io_x2 = m_453_io_cout; // @[MUL.scala 263:22]
  assign m_545_io_x3 = m_457_io_s; // @[MUL.scala 262:21]
  assign m_546_io_x1 = m_454_io_cout; // @[MUL.scala 263:22]
  assign m_546_io_x2 = m_158_io_cout; // @[MUL.scala 263:22]
  assign m_546_io_x3 = m_455_io_out_1; // @[MUL.scala 105:13]
  assign m_547_io_x1 = m_458_io_s; // @[MUL.scala 262:21]
  assign m_547_io_x2 = m_456_io_cout; // @[MUL.scala 263:22]
  assign m_547_io_x3 = m_459_io_s; // @[MUL.scala 262:21]
  assign m_548_io_in_0 = m_457_io_cout; // @[MUL.scala 263:22]
  assign m_548_io_in_1 = m_163_io_cout; // @[MUL.scala 263:22]
  assign m_549_io_x1 = m_460_io_s; // @[MUL.scala 262:21]
  assign m_549_io_x2 = m_458_io_cout; // @[MUL.scala 263:22]
  assign m_549_io_x3 = m_461_io_s; // @[MUL.scala 262:21]
  assign m_550_io_in_0 = m_459_io_cout; // @[MUL.scala 263:22]
  assign m_550_io_in_1 = m_168_io_out_1; // @[MUL.scala 126:16]
  assign m_551_io_x1 = m_462_io_s; // @[MUL.scala 262:21]
  assign m_551_io_x2 = m_460_io_cout; // @[MUL.scala 263:22]
  assign m_551_io_x3 = m_463_io_s; // @[MUL.scala 262:21]
  assign m_552_io_in_0 = m_461_io_cout; // @[MUL.scala 263:22]
  assign m_552_io_in_1 = m_173_io_out_1; // @[MUL.scala 126:16]
  assign m_553_io_x1 = m_464_io_s; // @[MUL.scala 262:21]
  assign m_553_io_x2 = m_462_io_cout; // @[MUL.scala 263:22]
  assign m_553_io_x3 = m_465_io_s; // @[MUL.scala 262:21]
  assign m_554_io_x1 = m_466_io_s; // @[MUL.scala 262:21]
  assign m_554_io_x2 = m_464_io_cout; // @[MUL.scala 263:22]
  assign m_554_io_x3 = m_467_io_s; // @[MUL.scala 262:21]
  assign m_555_io_x1 = m_468_io_s; // @[MUL.scala 262:21]
  assign m_555_io_x2 = m_466_io_cout; // @[MUL.scala 263:22]
  assign m_555_io_x3 = m_469_io_s; // @[MUL.scala 262:21]
  assign m_556_io_x1 = m_470_io_s; // @[MUL.scala 262:21]
  assign m_556_io_x2 = m_468_io_cout; // @[MUL.scala 263:22]
  assign m_556_io_x3 = m_471_io_s; // @[MUL.scala 262:21]
  assign m_557_io_x1 = m_472_io_s; // @[MUL.scala 262:21]
  assign m_557_io_x2 = m_470_io_cout; // @[MUL.scala 263:22]
  assign m_557_io_x3 = m_473_io_s; // @[MUL.scala 262:21]
  assign m_558_io_x1 = m_474_io_s; // @[MUL.scala 262:21]
  assign m_558_io_x2 = m_472_io_cout; // @[MUL.scala 263:22]
  assign m_558_io_x3 = m_475_io_s; // @[MUL.scala 262:21]
  assign m_559_io_x1 = m_476_io_s; // @[MUL.scala 262:21]
  assign m_559_io_x2 = m_474_io_cout; // @[MUL.scala 263:22]
  assign m_559_io_x3 = m_477_io_s; // @[MUL.scala 262:21]
  assign m_560_io_x1 = m_478_io_s; // @[MUL.scala 262:21]
  assign m_560_io_x2 = m_476_io_cout; // @[MUL.scala 263:22]
  assign m_560_io_x3 = m_362_io_cout; // @[MUL.scala 263:22]
  assign m_561_io_x1 = m_479_io_s; // @[MUL.scala 262:21]
  assign m_561_io_x2 = m_478_io_cout; // @[MUL.scala 263:22]
  assign m_561_io_x3 = m_364_io_cout; // @[MUL.scala 263:22]
  assign m_562_io_x1 = m_480_io_s; // @[MUL.scala 262:21]
  assign m_562_io_x2 = m_479_io_cout; // @[MUL.scala 263:22]
  assign m_562_io_x3 = m_366_io_cout; // @[MUL.scala 263:22]
  assign m_563_io_x1 = m_481_io_s; // @[MUL.scala 262:21]
  assign m_563_io_x2 = m_480_io_cout; // @[MUL.scala 263:22]
  assign m_563_io_x3 = m_368_io_cout; // @[MUL.scala 263:22]
  assign m_564_io_x1 = m_482_io_s; // @[MUL.scala 262:21]
  assign m_564_io_x2 = m_481_io_cout; // @[MUL.scala 263:22]
  assign m_564_io_x3 = m_370_io_cout; // @[MUL.scala 263:22]
  assign m_565_io_x1 = m_483_io_s; // @[MUL.scala 262:21]
  assign m_565_io_x2 = m_482_io_cout; // @[MUL.scala 263:22]
  assign m_565_io_x3 = m_372_io_cout; // @[MUL.scala 263:22]
  assign m_566_io_x1 = m_484_io_s; // @[MUL.scala 262:21]
  assign m_566_io_x2 = m_483_io_cout; // @[MUL.scala 263:22]
  assign m_566_io_x3 = m_374_io_out_1; // @[MUL.scala 105:13]
  assign m_567_io_in_0 = m_485_io_s; // @[MUL.scala 262:21]
  assign m_567_io_in_1 = m_484_io_cout; // @[MUL.scala 263:22]
  assign m_568_io_in_0 = m_486_io_s; // @[MUL.scala 262:21]
  assign m_568_io_in_1 = m_485_io_cout; // @[MUL.scala 263:22]
  assign m_569_io_in_0 = m_487_io_s; // @[MUL.scala 262:21]
  assign m_569_io_in_1 = m_486_io_cout; // @[MUL.scala 263:22]
  assign m_570_io_in_0 = m_488_io_s; // @[MUL.scala 262:21]
  assign m_570_io_in_1 = m_487_io_cout; // @[MUL.scala 263:22]
  assign m_571_io_in_0 = m_489_io_out_0; // @[MUL.scala 125:16]
  assign m_571_io_in_1 = m_488_io_cout; // @[MUL.scala 263:22]
  assign m_572_io_in_0 = m_490_io_out_0; // @[MUL.scala 125:16]
  assign m_572_io_in_1 = m_489_io_out_1; // @[MUL.scala 126:16]
  assign m_573_io_in_0 = m_491_io_out_0; // @[MUL.scala 125:16]
  assign m_573_io_in_1 = m_490_io_out_1; // @[MUL.scala 126:16]
  assign m_574_io_in_0 = m_492_io_out_0; // @[MUL.scala 125:16]
  assign m_574_io_in_1 = m_491_io_out_1; // @[MUL.scala 126:16]
  assign m_575_io_in_0 = m_493_io_out_0; // @[MUL.scala 125:16]
  assign m_575_io_in_1 = m_492_io_out_1; // @[MUL.scala 126:16]
  assign m_576_io_in_0 = m_494_io_out_0; // @[MUL.scala 125:16]
  assign m_576_io_in_1 = m_493_io_out_1; // @[MUL.scala 126:16]
  assign m_577_io_in_0 = r_648; // @[MUL.scala 125:16]
  assign m_577_io_in_1 = r_649; // @[MUL.scala 126:16]
  assign m_578_io_in_0 = r_650; // @[MUL.scala 125:16]
  assign m_578_io_in_1 = r_651; // @[MUL.scala 126:16]
  assign m_579_io_in_0 = r_652; // @[MUL.scala 125:16]
  assign m_579_io_in_1 = r_653; // @[MUL.scala 126:16]
  assign m_580_io_in_0 = r_654; // @[MUL.scala 125:16]
  assign m_580_io_in_1 = r_655; // @[MUL.scala 126:16]
  assign m_581_io_in_0 = r_656; // @[MUL.scala 125:16]
  assign m_581_io_in_1 = r_657; // @[MUL.scala 126:16]
  assign m_582_io_in_0 = r_658; // @[MUL.scala 125:16]
  assign m_582_io_in_1 = r_659; // @[MUL.scala 126:16]
  assign m_583_io_in_0 = r_660; // @[MUL.scala 125:16]
  assign m_583_io_in_1 = r_661; // @[MUL.scala 126:16]
  assign m_584_io_in_0 = r_662; // @[MUL.scala 125:16]
  assign m_584_io_in_1 = r_663; // @[MUL.scala 126:16]
  assign m_585_io_in_0 = r_664; // @[MUL.scala 125:16]
  assign m_585_io_in_1 = r_665; // @[MUL.scala 126:16]
  assign m_586_io_in_0 = r_666; // @[MUL.scala 125:16]
  assign m_586_io_in_1 = r_667; // @[MUL.scala 126:16]
  assign m_587_io_in_0 = r_668; // @[MUL.scala 125:16]
  assign m_587_io_in_1 = r_669; // @[MUL.scala 126:16]
  assign m_588_io_in_0 = r_670; // @[MUL.scala 125:16]
  assign m_588_io_in_1 = r_671; // @[MUL.scala 126:16]
  assign m_589_io_in_0 = r_672; // @[MUL.scala 125:16]
  assign m_589_io_in_1 = r_673; // @[MUL.scala 126:16]
  assign m_590_io_x1 = r_674; // @[MUL.scala 103:13]
  assign m_590_io_x2 = r_675; // @[MUL.scala 104:13]
  assign m_590_io_x3 = r_676; // @[MUL.scala 105:13]
  assign m_591_io_x1 = r_677; // @[MUL.scala 103:13]
  assign m_591_io_x2 = r_678; // @[MUL.scala 104:13]
  assign m_591_io_x3 = r_679; // @[MUL.scala 105:13]
  assign m_592_io_x1 = r_680; // @[MUL.scala 103:13]
  assign m_592_io_x2 = r_681; // @[MUL.scala 104:13]
  assign m_592_io_x3 = r_682; // @[MUL.scala 105:13]
  assign m_593_io_x1 = r_683; // @[MUL.scala 103:13]
  assign m_593_io_x2 = r_684; // @[MUL.scala 104:13]
  assign m_593_io_x3 = r_685; // @[MUL.scala 105:13]
  assign m_594_io_x1 = r_686; // @[MUL.scala 103:13]
  assign m_594_io_x2 = r_687; // @[MUL.scala 104:13]
  assign m_594_io_x3 = r_688; // @[MUL.scala 105:13]
  assign m_595_io_x1 = r_689; // @[MUL.scala 103:13]
  assign m_595_io_x2 = r_690; // @[MUL.scala 104:13]
  assign m_595_io_x3 = r_691; // @[MUL.scala 105:13]
  assign m_596_io_x1 = r_692; // @[MUL.scala 103:13]
  assign m_596_io_x2 = r_693; // @[MUL.scala 104:13]
  assign m_596_io_x3 = r_694; // @[MUL.scala 105:13]
  assign m_597_io_x1 = r_695; // @[MUL.scala 103:13]
  assign m_597_io_x2 = r_696; // @[MUL.scala 104:13]
  assign m_597_io_x3 = r_697; // @[MUL.scala 105:13]
  assign m_598_io_x1 = r_698; // @[MUL.scala 103:13]
  assign m_598_io_x2 = r_699; // @[MUL.scala 104:13]
  assign m_598_io_x3 = r_700; // @[MUL.scala 105:13]
  assign m_599_io_x1 = r_701; // @[MUL.scala 103:13]
  assign m_599_io_x2 = r_702; // @[MUL.scala 104:13]
  assign m_599_io_x3 = r_703; // @[MUL.scala 105:13]
  assign m_600_io_x1 = r_705; // @[MUL.scala 103:13]
  assign m_600_io_x2 = r_706; // @[MUL.scala 104:13]
  assign m_600_io_x3 = r_707; // @[MUL.scala 105:13]
  assign m_601_io_x1 = r_709; // @[MUL.scala 103:13]
  assign m_601_io_x2 = r_710; // @[MUL.scala 104:13]
  assign m_601_io_x3 = r_711; // @[MUL.scala 105:13]
  assign m_602_io_x1 = r_713; // @[MUL.scala 103:13]
  assign m_602_io_x2 = r_714; // @[MUL.scala 104:13]
  assign m_602_io_x3 = r_715; // @[MUL.scala 105:13]
  assign m_603_io_x1 = r_717; // @[MUL.scala 103:13]
  assign m_603_io_x2 = r_718; // @[MUL.scala 104:13]
  assign m_603_io_x3 = r_719; // @[MUL.scala 105:13]
  assign m_604_io_x1 = r_721; // @[MUL.scala 103:13]
  assign m_604_io_x2 = r_722; // @[MUL.scala 104:13]
  assign m_604_io_x3 = r_723; // @[MUL.scala 105:13]
  assign m_605_io_x1 = r_725; // @[MUL.scala 103:13]
  assign m_605_io_x2 = r_726; // @[MUL.scala 104:13]
  assign m_605_io_x3 = r_727; // @[MUL.scala 105:13]
  assign m_606_io_x1 = r_729; // @[MUL.scala 103:13]
  assign m_606_io_x2 = r_730; // @[MUL.scala 104:13]
  assign m_606_io_x3 = r_731; // @[MUL.scala 105:13]
  assign m_607_io_x1 = r_733; // @[MUL.scala 103:13]
  assign m_607_io_x2 = r_734; // @[MUL.scala 104:13]
  assign m_607_io_x3 = r_735; // @[MUL.scala 105:13]
  assign m_608_io_x1 = r_737; // @[MUL.scala 103:13]
  assign m_608_io_x2 = r_738; // @[MUL.scala 104:13]
  assign m_608_io_x3 = r_739; // @[MUL.scala 105:13]
  assign m_609_io_x1 = r_741; // @[MUL.scala 103:13]
  assign m_609_io_x2 = r_742; // @[MUL.scala 104:13]
  assign m_609_io_x3 = r_743; // @[MUL.scala 105:13]
  assign m_610_io_x1 = r_745; // @[MUL.scala 103:13]
  assign m_610_io_x2 = r_746; // @[MUL.scala 104:13]
  assign m_610_io_x3 = r_747; // @[MUL.scala 105:13]
  assign m_611_io_x1 = r_749; // @[MUL.scala 103:13]
  assign m_611_io_x2 = r_750; // @[MUL.scala 104:13]
  assign m_611_io_x3 = r_751; // @[MUL.scala 105:13]
  assign m_612_io_x1 = r_753; // @[MUL.scala 103:13]
  assign m_612_io_x2 = r_754; // @[MUL.scala 104:13]
  assign m_612_io_x3 = r_755; // @[MUL.scala 105:13]
  assign m_613_io_x1 = r_757; // @[MUL.scala 103:13]
  assign m_613_io_x2 = r_758; // @[MUL.scala 104:13]
  assign m_613_io_x3 = r_759; // @[MUL.scala 105:13]
  assign m_614_io_x1 = r_761; // @[MUL.scala 103:13]
  assign m_614_io_x2 = r_762; // @[MUL.scala 104:13]
  assign m_614_io_x3 = r_763; // @[MUL.scala 105:13]
  assign m_615_io_x1 = r_765; // @[MUL.scala 103:13]
  assign m_615_io_x2 = r_766; // @[MUL.scala 104:13]
  assign m_615_io_x3 = r_767; // @[MUL.scala 105:13]
  assign m_616_io_x1 = r_769; // @[MUL.scala 103:13]
  assign m_616_io_x2 = r_770; // @[MUL.scala 104:13]
  assign m_616_io_x3 = r_771; // @[MUL.scala 105:13]
  assign m_617_io_x1 = r_773; // @[MUL.scala 103:13]
  assign m_617_io_x2 = r_774; // @[MUL.scala 104:13]
  assign m_617_io_x3 = r_775; // @[MUL.scala 105:13]
  assign m_618_io_x1 = r_776; // @[MUL.scala 103:13]
  assign m_618_io_x2 = r_777; // @[MUL.scala 104:13]
  assign m_618_io_x3 = r_778; // @[MUL.scala 105:13]
  assign m_619_io_x1 = r_779; // @[MUL.scala 103:13]
  assign m_619_io_x2 = r_780; // @[MUL.scala 104:13]
  assign m_619_io_x3 = r_781; // @[MUL.scala 105:13]
  assign m_620_io_x1 = r_782; // @[MUL.scala 103:13]
  assign m_620_io_x2 = r_783; // @[MUL.scala 104:13]
  assign m_620_io_x3 = r_784; // @[MUL.scala 105:13]
  assign m_621_io_x1 = r_785; // @[MUL.scala 103:13]
  assign m_621_io_x2 = r_786; // @[MUL.scala 104:13]
  assign m_621_io_x3 = r_787; // @[MUL.scala 105:13]
  assign m_622_io_x1 = r_788; // @[MUL.scala 103:13]
  assign m_622_io_x2 = r_789; // @[MUL.scala 104:13]
  assign m_622_io_x3 = r_790; // @[MUL.scala 105:13]
  assign m_623_io_x1 = r_791; // @[MUL.scala 103:13]
  assign m_623_io_x2 = r_792; // @[MUL.scala 104:13]
  assign m_623_io_x3 = r_793; // @[MUL.scala 105:13]
  assign m_624_io_in_0 = r_794; // @[MUL.scala 125:16]
  assign m_624_io_in_1 = r_795; // @[MUL.scala 126:16]
  assign m_625_io_in_0 = r_796; // @[MUL.scala 125:16]
  assign m_625_io_in_1 = r_797; // @[MUL.scala 126:16]
  assign m_626_io_in_0 = r_798; // @[MUL.scala 125:16]
  assign m_626_io_in_1 = r_799; // @[MUL.scala 126:16]
  assign m_627_io_in_0 = r_800; // @[MUL.scala 125:16]
  assign m_627_io_in_1 = r_801; // @[MUL.scala 126:16]
  assign m_628_io_in_0 = r_802; // @[MUL.scala 125:16]
  assign m_628_io_in_1 = r_803; // @[MUL.scala 126:16]
  assign m_629_io_in_0 = r_804; // @[MUL.scala 125:16]
  assign m_629_io_in_1 = r_805; // @[MUL.scala 126:16]
  assign m_630_io_in_0 = r_806; // @[MUL.scala 125:16]
  assign m_630_io_in_1 = r_807; // @[MUL.scala 126:16]
  assign m_631_io_in_0 = r_808; // @[MUL.scala 125:16]
  assign m_631_io_in_1 = r_809; // @[MUL.scala 126:16]
  assign m_632_io_in_0 = r_810; // @[MUL.scala 125:16]
  assign m_632_io_in_1 = r_811; // @[MUL.scala 126:16]
  assign m_633_io_in_0 = r_812; // @[MUL.scala 125:16]
  assign m_633_io_in_1 = r_813; // @[MUL.scala 126:16]
  assign m_634_io_in_0 = r_814; // @[MUL.scala 125:16]
  assign m_634_io_in_1 = r_815; // @[MUL.scala 126:16]
  assign m_635_io_in_0 = r_816; // @[MUL.scala 125:16]
  assign m_635_io_in_1 = r_817; // @[MUL.scala 126:16]
  assign m_636_io_in_0 = r_818; // @[MUL.scala 125:16]
  assign m_636_io_in_1 = r_819; // @[MUL.scala 126:16]
  assign m_637_io_in_0 = r_820; // @[MUL.scala 125:16]
  assign m_637_io_in_1 = r_821; // @[MUL.scala 126:16]
  assign m_638_io_in_0 = r_822; // @[MUL.scala 125:16]
  assign m_638_io_in_1 = r_823; // @[MUL.scala 126:16]
  assign m_639_io_in_0 = r_824; // @[MUL.scala 125:16]
  assign m_639_io_in_1 = r_825; // @[MUL.scala 126:16]
  assign m_640_io_in_0 = m_578_io_out_0; // @[MUL.scala 125:16]
  assign m_640_io_in_1 = m_577_io_out_1; // @[MUL.scala 126:16]
  assign m_641_io_in_0 = m_579_io_out_0; // @[MUL.scala 125:16]
  assign m_641_io_in_1 = m_578_io_out_1; // @[MUL.scala 126:16]
  assign m_642_io_in_0 = m_580_io_out_0; // @[MUL.scala 125:16]
  assign m_642_io_in_1 = m_579_io_out_1; // @[MUL.scala 126:16]
  assign m_643_io_in_0 = m_581_io_out_0; // @[MUL.scala 125:16]
  assign m_643_io_in_1 = m_580_io_out_1; // @[MUL.scala 126:16]
  assign m_644_io_in_0 = m_582_io_out_0; // @[MUL.scala 125:16]
  assign m_644_io_in_1 = m_581_io_out_1; // @[MUL.scala 126:16]
  assign m_645_io_in_0 = m_583_io_out_0; // @[MUL.scala 125:16]
  assign m_645_io_in_1 = m_582_io_out_1; // @[MUL.scala 126:16]
  assign m_646_io_in_0 = m_584_io_out_0; // @[MUL.scala 125:16]
  assign m_646_io_in_1 = m_583_io_out_1; // @[MUL.scala 126:16]
  assign m_647_io_in_0 = m_585_io_out_0; // @[MUL.scala 125:16]
  assign m_647_io_in_1 = m_584_io_out_1; // @[MUL.scala 126:16]
  assign m_648_io_in_0 = m_586_io_out_0; // @[MUL.scala 125:16]
  assign m_648_io_in_1 = m_585_io_out_1; // @[MUL.scala 126:16]
  assign m_649_io_in_0 = m_587_io_out_0; // @[MUL.scala 125:16]
  assign m_649_io_in_1 = m_586_io_out_1; // @[MUL.scala 126:16]
  assign m_650_io_in_0 = m_588_io_out_0; // @[MUL.scala 125:16]
  assign m_650_io_in_1 = m_587_io_out_1; // @[MUL.scala 126:16]
  assign m_651_io_in_0 = m_589_io_out_0; // @[MUL.scala 125:16]
  assign m_651_io_in_1 = m_588_io_out_1; // @[MUL.scala 126:16]
  assign m_652_io_in_0 = m_590_io_s; // @[MUL.scala 262:21]
  assign m_652_io_in_1 = m_589_io_out_1; // @[MUL.scala 126:16]
  assign m_653_io_in_0 = m_591_io_s; // @[MUL.scala 262:21]
  assign m_653_io_in_1 = m_590_io_cout; // @[MUL.scala 263:22]
  assign m_654_io_in_0 = m_592_io_s; // @[MUL.scala 262:21]
  assign m_654_io_in_1 = m_591_io_cout; // @[MUL.scala 263:22]
  assign m_655_io_in_0 = m_593_io_s; // @[MUL.scala 262:21]
  assign m_655_io_in_1 = m_592_io_cout; // @[MUL.scala 263:22]
  assign m_656_io_in_0 = m_594_io_s; // @[MUL.scala 262:21]
  assign m_656_io_in_1 = m_593_io_cout; // @[MUL.scala 263:22]
  assign m_657_io_in_0 = m_595_io_s; // @[MUL.scala 262:21]
  assign m_657_io_in_1 = m_594_io_cout; // @[MUL.scala 263:22]
  assign m_658_io_in_0 = m_596_io_s; // @[MUL.scala 262:21]
  assign m_658_io_in_1 = m_595_io_cout; // @[MUL.scala 263:22]
  assign m_659_io_in_0 = m_597_io_s; // @[MUL.scala 262:21]
  assign m_659_io_in_1 = m_596_io_cout; // @[MUL.scala 263:22]
  assign m_660_io_in_0 = m_598_io_s; // @[MUL.scala 262:21]
  assign m_660_io_in_1 = m_597_io_cout; // @[MUL.scala 263:22]
  assign m_661_io_x1 = m_599_io_s; // @[MUL.scala 262:21]
  assign m_661_io_x2 = m_598_io_cout; // @[MUL.scala 263:22]
  assign m_661_io_x3 = r_704; // @[MUL.scala 105:13]
  assign m_662_io_x1 = m_600_io_s; // @[MUL.scala 262:21]
  assign m_662_io_x2 = m_599_io_cout; // @[MUL.scala 263:22]
  assign m_662_io_x3 = r_708; // @[MUL.scala 105:13]
  assign m_663_io_x1 = m_601_io_s; // @[MUL.scala 262:21]
  assign m_663_io_x2 = m_600_io_cout; // @[MUL.scala 263:22]
  assign m_663_io_x3 = r_712; // @[MUL.scala 105:13]
  assign m_664_io_x1 = m_602_io_s; // @[MUL.scala 262:21]
  assign m_664_io_x2 = m_601_io_cout; // @[MUL.scala 263:22]
  assign m_664_io_x3 = r_716; // @[MUL.scala 105:13]
  assign m_665_io_x1 = m_603_io_s; // @[MUL.scala 262:21]
  assign m_665_io_x2 = m_602_io_cout; // @[MUL.scala 263:22]
  assign m_665_io_x3 = r_720; // @[MUL.scala 105:13]
  assign m_666_io_x1 = m_604_io_s; // @[MUL.scala 262:21]
  assign m_666_io_x2 = m_603_io_cout; // @[MUL.scala 263:22]
  assign m_666_io_x3 = r_724; // @[MUL.scala 105:13]
  assign m_667_io_x1 = m_605_io_s; // @[MUL.scala 262:21]
  assign m_667_io_x2 = m_604_io_cout; // @[MUL.scala 263:22]
  assign m_667_io_x3 = r_728; // @[MUL.scala 105:13]
  assign m_668_io_x1 = m_606_io_s; // @[MUL.scala 262:21]
  assign m_668_io_x2 = m_605_io_cout; // @[MUL.scala 263:22]
  assign m_668_io_x3 = r_732; // @[MUL.scala 105:13]
  assign m_669_io_x1 = m_607_io_s; // @[MUL.scala 262:21]
  assign m_669_io_x2 = m_606_io_cout; // @[MUL.scala 263:22]
  assign m_669_io_x3 = r_736; // @[MUL.scala 105:13]
  assign m_670_io_x1 = m_608_io_s; // @[MUL.scala 262:21]
  assign m_670_io_x2 = m_607_io_cout; // @[MUL.scala 263:22]
  assign m_670_io_x3 = r_740; // @[MUL.scala 105:13]
  assign m_671_io_x1 = m_609_io_s; // @[MUL.scala 262:21]
  assign m_671_io_x2 = m_608_io_cout; // @[MUL.scala 263:22]
  assign m_671_io_x3 = r_744; // @[MUL.scala 105:13]
  assign m_672_io_x1 = m_610_io_s; // @[MUL.scala 262:21]
  assign m_672_io_x2 = m_609_io_cout; // @[MUL.scala 263:22]
  assign m_672_io_x3 = r_748; // @[MUL.scala 105:13]
  assign m_673_io_x1 = m_611_io_s; // @[MUL.scala 262:21]
  assign m_673_io_x2 = m_610_io_cout; // @[MUL.scala 263:22]
  assign m_673_io_x3 = r_752; // @[MUL.scala 105:13]
  assign m_674_io_x1 = m_612_io_s; // @[MUL.scala 262:21]
  assign m_674_io_x2 = m_611_io_cout; // @[MUL.scala 263:22]
  assign m_674_io_x3 = r_756; // @[MUL.scala 105:13]
  assign m_675_io_x1 = m_613_io_s; // @[MUL.scala 262:21]
  assign m_675_io_x2 = m_612_io_cout; // @[MUL.scala 263:22]
  assign m_675_io_x3 = r_760; // @[MUL.scala 105:13]
  assign m_676_io_x1 = m_614_io_s; // @[MUL.scala 262:21]
  assign m_676_io_x2 = m_613_io_cout; // @[MUL.scala 263:22]
  assign m_676_io_x3 = r_764; // @[MUL.scala 105:13]
  assign m_677_io_x1 = m_615_io_s; // @[MUL.scala 262:21]
  assign m_677_io_x2 = m_614_io_cout; // @[MUL.scala 263:22]
  assign m_677_io_x3 = r_768; // @[MUL.scala 105:13]
  assign m_678_io_x1 = m_616_io_s; // @[MUL.scala 262:21]
  assign m_678_io_x2 = m_615_io_cout; // @[MUL.scala 263:22]
  assign m_678_io_x3 = r_772; // @[MUL.scala 105:13]
  assign m_679_io_in_0 = m_617_io_s; // @[MUL.scala 262:21]
  assign m_679_io_in_1 = m_616_io_cout; // @[MUL.scala 263:22]
  assign m_680_io_in_0 = m_618_io_s; // @[MUL.scala 262:21]
  assign m_680_io_in_1 = m_617_io_cout; // @[MUL.scala 263:22]
  assign m_681_io_in_0 = m_619_io_s; // @[MUL.scala 262:21]
  assign m_681_io_in_1 = m_618_io_cout; // @[MUL.scala 263:22]
  assign m_682_io_in_0 = m_620_io_s; // @[MUL.scala 262:21]
  assign m_682_io_in_1 = m_619_io_cout; // @[MUL.scala 263:22]
  assign m_683_io_in_0 = m_621_io_s; // @[MUL.scala 262:21]
  assign m_683_io_in_1 = m_620_io_cout; // @[MUL.scala 263:22]
  assign m_684_io_in_0 = m_622_io_s; // @[MUL.scala 262:21]
  assign m_684_io_in_1 = m_621_io_cout; // @[MUL.scala 263:22]
  assign m_685_io_in_0 = m_623_io_s; // @[MUL.scala 262:21]
  assign m_685_io_in_1 = m_622_io_cout; // @[MUL.scala 263:22]
  assign m_686_io_in_0 = m_624_io_out_0; // @[MUL.scala 125:16]
  assign m_686_io_in_1 = m_623_io_cout; // @[MUL.scala 263:22]
  assign m_687_io_in_0 = m_625_io_out_0; // @[MUL.scala 125:16]
  assign m_687_io_in_1 = m_624_io_out_1; // @[MUL.scala 126:16]
  assign m_688_io_in_0 = m_626_io_out_0; // @[MUL.scala 125:16]
  assign m_688_io_in_1 = m_625_io_out_1; // @[MUL.scala 126:16]
  assign m_689_io_in_0 = m_627_io_out_0; // @[MUL.scala 125:16]
  assign m_689_io_in_1 = m_626_io_out_1; // @[MUL.scala 126:16]
  assign m_690_io_in_0 = m_628_io_out_0; // @[MUL.scala 125:16]
  assign m_690_io_in_1 = m_627_io_out_1; // @[MUL.scala 126:16]
  assign m_691_io_in_0 = m_629_io_out_0; // @[MUL.scala 125:16]
  assign m_691_io_in_1 = m_628_io_out_1; // @[MUL.scala 126:16]
  assign m_692_io_in_0 = m_630_io_out_0; // @[MUL.scala 125:16]
  assign m_692_io_in_1 = m_629_io_out_1; // @[MUL.scala 126:16]
  assign m_693_io_in_0 = m_631_io_out_0; // @[MUL.scala 125:16]
  assign m_693_io_in_1 = m_630_io_out_1; // @[MUL.scala 126:16]
  assign m_694_io_in_0 = m_632_io_out_0; // @[MUL.scala 125:16]
  assign m_694_io_in_1 = m_631_io_out_1; // @[MUL.scala 126:16]
  assign m_695_io_in_0 = m_633_io_out_0; // @[MUL.scala 125:16]
  assign m_695_io_in_1 = m_632_io_out_1; // @[MUL.scala 126:16]
  assign m_696_io_in_0 = m_634_io_out_0; // @[MUL.scala 125:16]
  assign m_696_io_in_1 = m_633_io_out_1; // @[MUL.scala 126:16]
  assign m_697_io_in_0 = m_635_io_out_0; // @[MUL.scala 125:16]
  assign m_697_io_in_1 = m_634_io_out_1; // @[MUL.scala 126:16]
  assign m_698_io_in_0 = m_636_io_out_0; // @[MUL.scala 125:16]
  assign m_698_io_in_1 = m_635_io_out_1; // @[MUL.scala 126:16]
  assign m_699_io_in_0 = m_637_io_out_0; // @[MUL.scala 125:16]
  assign m_699_io_in_1 = m_636_io_out_1; // @[MUL.scala 126:16]
  assign m_700_io_in_0 = m_638_io_out_0; // @[MUL.scala 125:16]
  assign m_700_io_in_1 = m_637_io_out_1; // @[MUL.scala 126:16]
  assign m_701_io_in_0 = m_639_io_out_0; // @[MUL.scala 125:16]
  assign m_701_io_in_1 = m_638_io_out_1; // @[MUL.scala 126:16]
  always @(posedge clock) begin
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r <= m_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_1 <= m_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_2 <= m_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_3 <= m_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_4 <= m_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_5 <= m_1_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_6 <= m_1_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_7 <= m_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_8 <= m_1_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_9 <= m_1_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_10 <= m_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_11 <= m_1_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_12 <= m_2_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_13 <= m_2_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_14 <= m_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_15 <= m_1_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_16 <= m_2_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_17 <= m_2_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_18 <= m_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_19 <= m_1_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_20 <= m_2_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_21 <= m_3_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_22 <= m_3_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_23 <= m_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_24 <= m_1_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_25 <= m_2_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_26 <= m_3_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_27 <= m_3_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_28 <= m_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_29 <= m_1_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_30 <= m_2_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_31 <= m_3_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_32 <= m_4_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_33 <= m_4_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_34 <= m_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_35 <= m_1_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_36 <= m_2_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_37 <= m_3_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_38 <= m_4_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_39 <= m_4_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_40 <= m_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_41 <= m_1_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_42 <= m_2_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_43 <= m_3_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_44 <= m_4_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_45 <= m_5_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_46 <= m_5_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_47 <= m_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_48 <= m_1_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_49 <= m_2_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_50 <= m_3_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_51 <= m_4_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_52 <= m_5_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_53 <= m_5_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_54 <= m_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_55 <= m_1_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_56 <= m_2_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_57 <= m_3_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_58 <= m_4_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_59 <= m_5_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_60 <= m_6_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_61 <= m_6_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_62 <= m_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_63 <= m_1_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_64 <= m_2_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_65 <= m_3_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_66 <= m_4_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_67 <= m_5_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_68 <= m_6_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_69 <= m_6_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_70 <= m_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_71 <= m_1_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_72 <= m_2_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_73 <= m_3_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_74 <= m_4_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_75 <= m_5_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_76 <= m_6_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_77 <= m_7_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_78 <= m_7_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_79 <= m_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_80 <= m_1_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_81 <= m_2_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_82 <= m_3_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_83 <= m_4_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_84 <= m_5_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_85 <= m_6_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_86 <= m_7_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_87 <= m_7_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_88 <= m_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_89 <= m_1_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_90 <= m_2_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_91 <= m_3_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_92 <= m_4_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_93 <= m_5_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_94 <= m_6_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_95 <= m_7_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_96 <= m_8_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_97 <= m_8_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_98 <= m_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_99 <= m_1_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_100 <= m_2_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_101 <= m_3_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_102 <= m_4_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_103 <= m_5_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_104 <= m_6_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_105 <= m_7_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_106 <= m_8_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_107 <= m_8_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_108 <= m_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_109 <= m_1_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_110 <= m_2_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_111 <= m_3_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_112 <= m_4_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_113 <= m_5_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_114 <= m_6_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_115 <= m_7_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_116 <= m_8_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_117 <= m_9_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_118 <= m_9_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_119 <= m_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_120 <= m_1_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_121 <= m_2_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_122 <= m_3_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_123 <= m_4_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_124 <= m_5_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_125 <= m_6_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_126 <= m_7_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_127 <= m_8_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_128 <= m_9_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_129 <= m_9_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_130 <= m_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_131 <= m_1_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_132 <= m_2_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_133 <= m_3_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_134 <= m_4_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_135 <= m_5_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_136 <= m_6_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_137 <= m_7_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_138 <= m_8_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_139 <= m_9_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_140 <= m_10_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_141 <= m_10_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_142 <= m_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_143 <= m_1_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_144 <= m_2_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_145 <= m_3_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_146 <= m_4_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_147 <= m_5_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_148 <= m_6_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_149 <= m_7_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_150 <= m_8_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_151 <= m_9_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_152 <= m_10_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_153 <= m_10_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_154 <= m_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_155 <= m_1_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_156 <= m_2_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_157 <= m_3_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_158 <= m_4_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_159 <= m_5_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_160 <= m_6_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_161 <= m_7_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_162 <= m_8_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_163 <= m_9_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_164 <= m_10_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_165 <= m_11_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_166 <= m_11_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_167 <= m_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_168 <= m_1_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_169 <= m_2_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_170 <= m_3_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_171 <= m_4_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_172 <= m_5_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_173 <= m_6_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_174 <= m_7_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_175 <= m_8_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_176 <= m_9_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_177 <= m_10_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_178 <= m_11_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_179 <= m_11_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_180 <= m_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_181 <= m_1_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_182 <= m_2_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_183 <= m_3_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_184 <= m_4_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_185 <= m_5_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_186 <= m_6_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_187 <= m_7_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_188 <= m_8_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_189 <= m_9_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_190 <= m_10_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_191 <= m_11_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_192 <= m_12_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_193 <= m_12_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_194 <= m_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_195 <= m_1_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_196 <= m_2_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_197 <= m_3_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_198 <= m_4_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_199 <= m_5_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_200 <= m_6_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_201 <= m_7_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_202 <= m_8_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_203 <= m_9_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_204 <= m_10_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_205 <= m_11_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_206 <= m_12_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_207 <= m_12_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_208 <= m_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_209 <= m_1_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_210 <= m_2_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_211 <= m_3_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_212 <= m_4_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_213 <= m_5_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_214 <= m_6_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_215 <= m_7_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_216 <= m_8_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_217 <= m_9_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_218 <= m_10_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_219 <= m_11_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_220 <= m_12_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_221 <= m_13_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_222 <= m_13_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_223 <= m_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_224 <= m_1_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_225 <= m_2_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_226 <= m_3_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_227 <= m_4_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_228 <= m_5_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_229 <= m_6_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_230 <= m_7_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_231 <= m_8_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_232 <= m_9_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_233 <= m_10_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_234 <= m_11_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_235 <= m_12_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_236 <= m_13_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_237 <= m_13_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_238 <= m_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_239 <= m_1_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_240 <= m_2_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_241 <= m_3_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_242 <= m_4_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_243 <= m_5_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_244 <= m_6_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_245 <= m_7_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_246 <= m_8_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_247 <= m_9_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_248 <= m_10_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_249 <= m_11_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_250 <= m_12_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_251 <= m_13_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_252 <= m_14_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_253 <= m_14_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_254 <= m_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_255 <= m_1_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_256 <= m_2_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_257 <= m_3_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_258 <= m_4_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_259 <= m_5_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_260 <= m_6_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_261 <= m_7_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_262 <= m_8_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_263 <= m_9_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_264 <= m_10_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_265 <= m_11_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_266 <= m_12_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_267 <= m_13_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_268 <= m_14_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_269 <= m_14_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_270 <= m_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_271 <= m_1_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_272 <= m_2_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_273 <= m_3_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_274 <= m_4_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_275 <= m_5_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_276 <= m_6_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_277 <= m_7_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_278 <= m_8_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_279 <= m_9_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_280 <= m_10_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_281 <= m_11_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_282 <= m_12_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_283 <= m_13_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_284 <= m_14_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_285 <= m_15_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_286 <= m_15_io_carry[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_287 <= m_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_288 <= m_1_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_289 <= m_2_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_290 <= m_3_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_291 <= m_4_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_292 <= m_5_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_293 <= m_6_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_294 <= m_7_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_295 <= m_8_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_296 <= m_9_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_297 <= m_10_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_298 <= m_11_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_299 <= m_12_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_300 <= m_13_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_301 <= m_14_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_302 <= m_15_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_303 <= m_15_io_carry[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_304 <= m_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_305 <= m_1_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_306 <= m_2_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_307 <= m_3_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_308 <= m_4_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_309 <= m_5_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_310 <= m_6_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_311 <= m_7_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_312 <= m_8_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_313 <= m_9_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_314 <= m_10_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_315 <= m_11_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_316 <= m_12_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_317 <= m_13_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_318 <= m_14_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_319 <= m_15_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_320 <= m_16_io_p[0]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_321 <= m_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_322 <= m_1_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_323 <= m_2_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_324 <= m_3_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_325 <= m_4_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_326 <= m_5_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_327 <= m_6_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_328 <= m_7_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_329 <= m_8_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_330 <= m_9_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_331 <= m_10_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_332 <= m_11_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_333 <= m_12_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_334 <= m_13_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_335 <= m_14_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_336 <= m_15_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_337 <= m_16_io_p[1]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_338 <= m_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_339 <= m_1_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_340 <= m_2_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_341 <= m_3_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_342 <= m_4_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_343 <= m_5_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_344 <= m_6_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_345 <= m_7_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_346 <= m_8_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_347 <= m_9_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_348 <= m_10_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_349 <= m_11_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_350 <= m_12_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_351 <= m_13_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_352 <= m_14_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_353 <= m_15_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_354 <= m_16_io_p[2]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_355 <= m_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_356 <= m_1_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_357 <= m_2_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_358 <= m_3_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_359 <= m_4_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_360 <= m_5_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_361 <= m_6_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_362 <= m_7_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_363 <= m_8_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_364 <= m_9_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_365 <= m_10_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_366 <= m_11_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_367 <= m_12_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_368 <= m_13_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_369 <= m_14_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_370 <= m_15_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_371 <= m_16_io_p[3]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_372 <= _T_56; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_373 <= _T_93; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_374 <= m_2_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_375 <= m_3_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_376 <= m_4_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_377 <= m_5_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_378 <= m_6_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_379 <= m_7_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_380 <= m_8_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_381 <= m_9_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_382 <= m_10_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_383 <= m_11_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_384 <= m_12_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_385 <= m_13_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_386 <= m_14_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_387 <= m_15_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_388 <= m_16_io_p[4]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_390 <= m_2_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_391 <= m_3_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_392 <= m_4_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_393 <= m_5_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_394 <= m_6_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_395 <= m_7_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_396 <= m_8_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_397 <= m_9_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_398 <= m_10_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_399 <= m_11_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_400 <= m_12_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_401 <= m_13_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_402 <= m_14_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_403 <= m_15_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_404 <= m_16_io_p[5]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_405 <= _T_132; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_406 <= m_3_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_407 <= m_4_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_408 <= m_5_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_409 <= m_6_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_410 <= m_7_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_411 <= m_8_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_412 <= m_9_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_413 <= m_10_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_414 <= m_11_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_415 <= m_12_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_416 <= m_13_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_417 <= m_14_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_418 <= m_15_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_419 <= m_16_io_p[6]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_421 <= m_3_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_422 <= m_4_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_423 <= m_5_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_424 <= m_6_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_425 <= m_7_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_426 <= m_8_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_427 <= m_9_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_428 <= m_10_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_429 <= m_11_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_430 <= m_12_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_431 <= m_13_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_432 <= m_14_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_433 <= m_15_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_434 <= m_16_io_p[7]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_435 <= _T_171; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_436 <= m_4_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_437 <= m_5_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_438 <= m_6_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_439 <= m_7_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_440 <= m_8_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_441 <= m_9_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_442 <= m_10_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_443 <= m_11_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_444 <= m_12_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_445 <= m_13_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_446 <= m_14_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_447 <= m_15_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_448 <= m_16_io_p[8]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_450 <= m_4_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_451 <= m_5_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_452 <= m_6_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_453 <= m_7_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_454 <= m_8_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_455 <= m_9_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_456 <= m_10_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_457 <= m_11_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_458 <= m_12_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_459 <= m_13_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_460 <= m_14_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_461 <= m_15_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_462 <= m_16_io_p[9]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_463 <= _T_210; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_464 <= m_5_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_465 <= m_6_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_466 <= m_7_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_467 <= m_8_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_468 <= m_9_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_469 <= m_10_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_470 <= m_11_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_471 <= m_12_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_472 <= m_13_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_473 <= m_14_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_474 <= m_15_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_475 <= m_16_io_p[10]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_477 <= m_5_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_478 <= m_6_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_479 <= m_7_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_480 <= m_8_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_481 <= m_9_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_482 <= m_10_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_483 <= m_11_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_484 <= m_12_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_485 <= m_13_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_486 <= m_14_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_487 <= m_15_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_488 <= m_16_io_p[11]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_489 <= _T_249; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_490 <= m_6_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_491 <= m_7_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_492 <= m_8_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_493 <= m_9_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_494 <= m_10_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_495 <= m_11_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_496 <= m_12_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_497 <= m_13_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_498 <= m_14_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_499 <= m_15_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_500 <= m_16_io_p[12]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_502 <= m_6_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_503 <= m_7_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_504 <= m_8_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_505 <= m_9_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_506 <= m_10_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_507 <= m_11_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_508 <= m_12_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_509 <= m_13_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_510 <= m_14_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_511 <= m_15_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_512 <= m_16_io_p[13]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_513 <= _T_288; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_514 <= m_7_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_515 <= m_8_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_516 <= m_9_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_517 <= m_10_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_518 <= m_11_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_519 <= m_12_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_520 <= m_13_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_521 <= m_14_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_522 <= m_15_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_523 <= m_16_io_p[14]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_525 <= m_7_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_526 <= m_8_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_527 <= m_9_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_528 <= m_10_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_529 <= m_11_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_530 <= m_12_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_531 <= m_13_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_532 <= m_14_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_533 <= m_15_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_534 <= m_16_io_p[15]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_535 <= _T_327; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_536 <= m_8_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_537 <= m_9_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_538 <= m_10_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_539 <= m_11_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_540 <= m_12_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_541 <= m_13_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_542 <= m_14_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_543 <= m_15_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_544 <= m_16_io_p[16]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_546 <= m_8_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_547 <= m_9_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_548 <= m_10_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_549 <= m_11_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_550 <= m_12_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_551 <= m_13_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_552 <= m_14_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_553 <= m_15_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_554 <= m_16_io_p[17]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_555 <= _T_366; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_556 <= m_9_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_557 <= m_10_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_558 <= m_11_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_559 <= m_12_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_560 <= m_13_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_561 <= m_14_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_562 <= m_15_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_563 <= m_16_io_p[18]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_565 <= m_9_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_566 <= m_10_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_567 <= m_11_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_568 <= m_12_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_569 <= m_13_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_570 <= m_14_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_571 <= m_15_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_572 <= m_16_io_p[19]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_573 <= _T_405; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_574 <= m_10_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_575 <= m_11_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_576 <= m_12_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_577 <= m_13_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_578 <= m_14_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_579 <= m_15_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_580 <= m_16_io_p[20]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_582 <= m_10_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_583 <= m_11_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_584 <= m_12_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_585 <= m_13_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_586 <= m_14_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_587 <= m_15_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_588 <= m_16_io_p[21]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_589 <= _T_444; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_590 <= m_11_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_591 <= m_12_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_592 <= m_13_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_593 <= m_14_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_594 <= m_15_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_595 <= m_16_io_p[22]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_597 <= m_11_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_598 <= m_12_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_599 <= m_13_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_600 <= m_14_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_601 <= m_15_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_602 <= m_16_io_p[23]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_603 <= _T_483; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_604 <= m_12_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_605 <= m_13_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_606 <= m_14_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_607 <= m_15_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_608 <= m_16_io_p[24]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_610 <= m_12_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_611 <= m_13_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_612 <= m_14_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_613 <= m_15_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_614 <= m_16_io_p[25]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_615 <= _T_522; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_616 <= m_13_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_617 <= m_14_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_618 <= m_15_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_619 <= m_16_io_p[26]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_621 <= m_13_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_622 <= m_14_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_623 <= m_15_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_624 <= m_16_io_p[27]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_625 <= _T_561; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_626 <= m_14_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_627 <= m_15_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_628 <= m_16_io_p[28]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_630 <= m_14_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_631 <= m_15_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_632 <= m_16_io_p[29]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_633 <= _T_600; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_634 <= m_15_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_635 <= m_16_io_p[30]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_637 <= m_15_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_638 <= m_16_io_p[31]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_639 <= _T_639; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_640 <= m_16_io_p[32]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_642 <= m_16_io_p[33]; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_643 <= _T_678; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_644 <= m_17_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_645 <= m_234_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_646 <= m_386_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_647 <= m_495_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_648 <= m_496_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_649 <= m_495_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_650 <= m_497_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_651 <= m_496_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_652 <= m_498_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_653 <= m_497_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_654 <= m_499_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_655 <= m_498_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_656 <= m_500_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_657 <= m_499_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_658 <= m_501_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_659 <= m_500_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_660 <= m_502_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_661 <= m_501_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_662 <= s_0_174; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_663 <= m_502_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_664 <= s_0_175; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_665 <= c_0_174; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_666 <= s_0_176; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_667 <= c_0_175; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_668 <= s_0_177; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_669 <= c_0_176; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_670 <= s_0_178; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_671 <= c_0_177; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_672 <= s_0_179; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_673 <= c_0_178; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_674 <= s_0_180; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_675 <= c_0_179; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_676 <= m_401_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_677 <= s_0_181; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_678 <= c_0_180; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_679 <= m_403_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_680 <= s_0_182; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_681 <= c_0_181; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_682 <= m_405_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_683 <= s_0_183; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_684 <= c_0_182; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_685 <= m_407_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_686 <= s_0_184; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_687 <= c_0_183; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_688 <= c_1_92; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_689 <= s_0_185; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_690 <= c_0_184; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_691 <= c_1_93; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_692 <= s_0_186; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_693 <= c_0_185; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_694 <= c_1_94; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_695 <= s_0_187; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_696 <= c_0_186; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_697 <= c_1_95; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_698 <= s_0_188; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_699 <= c_0_187; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_700 <= m_518_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_701 <= s_0_189; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_702 <= c_0_188; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_703 <= m_520_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_704 <= m_518_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_705 <= s_0_190; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_706 <= c_0_189; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_707 <= m_522_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_708 <= m_520_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_709 <= s_0_191; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_710 <= c_0_190; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_711 <= m_524_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_712 <= m_522_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_713 <= s_0_192; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_714 <= c_0_191; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_715 <= m_526_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_716 <= m_524_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_717 <= s_0_193; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_718 <= c_0_192; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_719 <= s_2_122; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_720 <= m_526_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_721 <= s_0_194; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_722 <= c_0_193; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_723 <= s_2_123; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_724 <= c_1_122; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_725 <= s_0_195; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_726 <= c_0_194; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_727 <= s_2_124; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_728 <= c_1_123; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_729 <= s_0_196; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_730 <= c_0_195; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_731 <= s_2_125; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_732 <= c_1_124; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_733 <= s_0_197; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_734 <= c_0_196; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_735 <= s_2_126; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_736 <= c_1_125; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_737 <= s_0_198; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_738 <= c_0_197; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_739 <= s_2_127; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_740 <= c_1_126; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_741 <= s_0_199; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_742 <= c_0_198; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_743 <= s_2_128; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_744 <= c_1_127; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_745 <= s_0_200; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_746 <= c_0_199; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_747 <= s_2_129; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_748 <= c_1_128; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_749 <= s_0_201; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_750 <= c_0_200; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_751 <= s_2_130; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_752 <= c_1_129; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_753 <= s_0_202; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_754 <= c_0_201; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_755 <= s_2_131; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_756 <= c_1_130; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_757 <= s_0_203; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_758 <= c_0_202; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_759 <= m_548_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_760 <= c_1_131; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_761 <= s_0_204; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_762 <= c_0_203; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_763 <= m_550_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_764 <= m_548_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_765 <= s_0_205; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_766 <= c_0_204; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_767 <= m_552_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_768 <= m_550_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_769 <= s_0_206; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_770 <= c_0_205; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_771 <= c_1_114; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_772 <= m_552_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_773 <= s_0_207; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_774 <= c_0_206; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_775 <= c_1_115; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_776 <= s_0_208; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_777 <= c_0_207; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_778 <= c_1_116; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_779 <= s_0_209; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_780 <= c_0_208; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_781 <= c_1_117; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_782 <= s_0_210; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_783 <= c_0_209; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_784 <= c_1_118; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_785 <= s_0_211; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_786 <= c_0_210; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_787 <= c_1_119; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_788 <= s_0_212; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_789 <= c_0_211; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_790 <= c_1_120; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_791 <= s_0_213; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_792 <= c_0_212; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_793 <= c_1_121; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_794 <= s_0_214; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_795 <= c_0_213; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_796 <= s_0_215; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_797 <= c_0_214; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_798 <= s_0_216; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_799 <= c_0_215; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_800 <= s_0_217; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_801 <= c_0_216; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_802 <= s_0_218; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_803 <= c_0_217; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_804 <= s_0_219; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_805 <= c_0_218; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_806 <= m_567_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_807 <= c_0_219; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_808 <= m_568_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_809 <= m_567_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_810 <= m_569_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_811 <= m_568_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_812 <= m_570_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_813 <= m_569_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_814 <= m_571_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_815 <= m_570_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_816 <= m_572_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_817 <= m_571_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_818 <= m_573_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_819 <= m_572_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_820 <= m_574_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_821 <= m_573_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_822 <= m_575_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_823 <= m_574_io_out_1; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_824 <= m_576_io_out_0; // @[Reg.scala 20:22]
    end
    if (io_in_valid) begin // @[Reg.scala 20:18]
      r_825 <= m_575_io_out_1; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[MUL.scala 344:22]
      count <= 8'h0; // @[MUL.scala 344:22]
    end else if (~io_in_bits_ctrl_flow_flush & io_in_valid & ~io_out_valid) begin // @[MUL.scala 346:15]
      count <= _count_T_5;
    end else begin
      count <= 8'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  r_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  r_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  r_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  r_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  r_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  r_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  r_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  r_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  r_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  r_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  r_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  r_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  r_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  r_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  r_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  r_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  r_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  r_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  r_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  r_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  r_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  r_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  r_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  r_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  r_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  r_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  r_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  r_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  r_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  r_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  r_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  r_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  r_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  r_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  r_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  r_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  r_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  r_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  r_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  r_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  r_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  r_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  r_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  r_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  r_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  r_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  r_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  r_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  r_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  r_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  r_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  r_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  r_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  r_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  r_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  r_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  r_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  r_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  r_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  r_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  r_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  r_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  r_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  r_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  r_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  r_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  r_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  r_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  r_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  r_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  r_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  r_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  r_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  r_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  r_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  r_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  r_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  r_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  r_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  r_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  r_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  r_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  r_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  r_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  r_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  r_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  r_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  r_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  r_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  r_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  r_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  r_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  r_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  r_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  r_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  r_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  r_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  r_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  r_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  r_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  r_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  r_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  r_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  r_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  r_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  r_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  r_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  r_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  r_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  r_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  r_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  r_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  r_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  r_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  r_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  r_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  r_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  r_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  r_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  r_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  r_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  r_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  r_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  r_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  r_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  r_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  r_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  r_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  r_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  r_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  r_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  r_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  r_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  r_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  r_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  r_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  r_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  r_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  r_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  r_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  r_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  r_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  r_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  r_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  r_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  r_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  r_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  r_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  r_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  r_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  r_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  r_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  r_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  r_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  r_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  r_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  r_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  r_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  r_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  r_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  r_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  r_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  r_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  r_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  r_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  r_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  r_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  r_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  r_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  r_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  r_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  r_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  r_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  r_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  r_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  r_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  r_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  r_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  r_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  r_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  r_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  r_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  r_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  r_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  r_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  r_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  r_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  r_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  r_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  r_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  r_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  r_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  r_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  r_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  r_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  r_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  r_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  r_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  r_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  r_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  r_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  r_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  r_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  r_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  r_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  r_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  r_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  r_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  r_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  r_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  r_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  r_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  r_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  r_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  r_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  r_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  r_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  r_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  r_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  r_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  r_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  r_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  r_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  r_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  r_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  r_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  r_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  r_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  r_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  r_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  r_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  r_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  r_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  r_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  r_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  r_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  r_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  r_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  r_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  r_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  r_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  r_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  r_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  r_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  r_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  r_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  r_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  r_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  r_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  r_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  r_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  r_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  r_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  r_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  r_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  r_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  r_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  r_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  r_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  r_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  r_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  r_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  r_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  r_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  r_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  r_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  r_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  r_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  r_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  r_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  r_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  r_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  r_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  r_390 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  r_391 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  r_392 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  r_393 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  r_394 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  r_395 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  r_396 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  r_397 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  r_398 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  r_399 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  r_400 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  r_401 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  r_402 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  r_403 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  r_404 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  r_405 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  r_406 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  r_407 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  r_408 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  r_409 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  r_410 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  r_411 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  r_412 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  r_413 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  r_414 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  r_415 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  r_416 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  r_417 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  r_418 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  r_419 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  r_421 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  r_422 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  r_423 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  r_424 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  r_425 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  r_426 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  r_427 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  r_428 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  r_429 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  r_430 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  r_431 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  r_432 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  r_433 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  r_434 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  r_435 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  r_436 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  r_437 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  r_438 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  r_439 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  r_440 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  r_441 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  r_442 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  r_443 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  r_444 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  r_445 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  r_446 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  r_447 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  r_448 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  r_450 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  r_451 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  r_452 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  r_453 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  r_454 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  r_455 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  r_456 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  r_457 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  r_458 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  r_459 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  r_460 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  r_461 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  r_462 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  r_463 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  r_464 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  r_465 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  r_466 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  r_467 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  r_468 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  r_469 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  r_470 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  r_471 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  r_472 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  r_473 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  r_474 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  r_475 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  r_477 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  r_478 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  r_479 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  r_480 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  r_481 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  r_482 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  r_483 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  r_484 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  r_485 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  r_486 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  r_487 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  r_488 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  r_489 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  r_490 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  r_491 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  r_492 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  r_493 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  r_494 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  r_495 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  r_496 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  r_497 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  r_498 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  r_499 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  r_500 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  r_502 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  r_503 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  r_504 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  r_505 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  r_506 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  r_507 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  r_508 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  r_509 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  r_510 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  r_511 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  r_512 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  r_513 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  r_514 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  r_515 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  r_516 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  r_517 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  r_518 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  r_519 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  r_520 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  r_521 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  r_522 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  r_523 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  r_525 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  r_526 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  r_527 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  r_528 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  r_529 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  r_530 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  r_531 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  r_532 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  r_533 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  r_534 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  r_535 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  r_536 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  r_537 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  r_538 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  r_539 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  r_540 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  r_541 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  r_542 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  r_543 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  r_544 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  r_546 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  r_547 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  r_548 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  r_549 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  r_550 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  r_551 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  r_552 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  r_553 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  r_554 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  r_555 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  r_556 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  r_557 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  r_558 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  r_559 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  r_560 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  r_561 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  r_562 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  r_563 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  r_565 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  r_566 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  r_567 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  r_568 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  r_569 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  r_570 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  r_571 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  r_572 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  r_573 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  r_574 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  r_575 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  r_576 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  r_577 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  r_578 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  r_579 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  r_580 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  r_582 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  r_583 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  r_584 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  r_585 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  r_586 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  r_587 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  r_588 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  r_589 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  r_590 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  r_591 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  r_592 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  r_593 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  r_594 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  r_595 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  r_597 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  r_598 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  r_599 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  r_600 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  r_601 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  r_602 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  r_603 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  r_604 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  r_605 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  r_606 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  r_607 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  r_608 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  r_610 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  r_611 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  r_612 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  r_613 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  r_614 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  r_615 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  r_616 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  r_617 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  r_618 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  r_619 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  r_621 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  r_622 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  r_623 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  r_624 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  r_625 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  r_626 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  r_627 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  r_628 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  r_630 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  r_631 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  r_632 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  r_633 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  r_634 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  r_635 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  r_637 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  r_638 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  r_639 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  r_640 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  r_642 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  r_643 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  r_644 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  r_645 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  r_646 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  r_647 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  r_648 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  r_649 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  r_650 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  r_651 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  r_652 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  r_653 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  r_654 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  r_655 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  r_656 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  r_657 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  r_658 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  r_659 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  r_660 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  r_661 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  r_662 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  r_663 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  r_664 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  r_665 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  r_666 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  r_667 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  r_668 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  r_669 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  r_670 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  r_671 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  r_672 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  r_673 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  r_674 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  r_675 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  r_676 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  r_677 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  r_678 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  r_679 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  r_680 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  r_681 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  r_682 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  r_683 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  r_684 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  r_685 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  r_686 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  r_687 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  r_688 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  r_689 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  r_690 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  r_691 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  r_692 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  r_693 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  r_694 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  r_695 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  r_696 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  r_697 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  r_698 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  r_699 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  r_700 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  r_701 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  r_702 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  r_703 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  r_704 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  r_705 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  r_706 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  r_707 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  r_708 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  r_709 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  r_710 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  r_711 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  r_712 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  r_713 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  r_714 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  r_715 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  r_716 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  r_717 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  r_718 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  r_719 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  r_720 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  r_721 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  r_722 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  r_723 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  r_724 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  r_725 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  r_726 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  r_727 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  r_728 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  r_729 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  r_730 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  r_731 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  r_732 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  r_733 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  r_734 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  r_735 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  r_736 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  r_737 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  r_738 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  r_739 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  r_740 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  r_741 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  r_742 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  r_743 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  r_744 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  r_745 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  r_746 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  r_747 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  r_748 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  r_749 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  r_750 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  r_751 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  r_752 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  r_753 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  r_754 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  r_755 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  r_756 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  r_757 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  r_758 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  r_759 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  r_760 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  r_761 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  r_762 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  r_763 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  r_764 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  r_765 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  r_766 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  r_767 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  r_768 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  r_769 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  r_770 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  r_771 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  r_772 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  r_773 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  r_774 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  r_775 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  r_776 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  r_777 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  r_778 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  r_779 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  r_780 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  r_781 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  r_782 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  r_783 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  r_784 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  r_785 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  r_786 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  r_787 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  r_788 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  r_789 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  r_790 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  r_791 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  r_792 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  r_793 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  r_794 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  r_795 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  r_796 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  r_797 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  r_798 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  r_799 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  r_800 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  r_801 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  r_802 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  r_803 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  r_804 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  r_805 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  r_806 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  r_807 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  r_808 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  r_809 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  r_810 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  r_811 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  r_812 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  r_813 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  r_814 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  r_815 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  r_816 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  r_817 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  r_818 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  r_819 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  r_820 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  r_821 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  r_822 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  r_823 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  r_824 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  r_825 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  count = _RAND_811[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule


