
module ID (
    input [31:0] Inst//inst from inst ram
    output [7:0] InstOP,
    output [3:0] InstType,
    output [2:0] ALUop
);





endmodule //ID