`define RestEn 1'b1
`define RestDis 1'b0
`define false 1'b0
`define true 1'b1
`define bypass_width 38
`define ctrl_width 211
`define ex_ctrl_width 220
`define mem_ctrl_width 104