
module ID (
    input [31:0] Inst//inst from inst ram
    output []
);





endmodule //ID