
module Top (
    ports
);
    
endmodule

